

package multi_queue_fifo_reader_pkg;

endpackage

interface multi_queue_fifo_reader_out_stream_if import multi_queue_fifo_reader_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface multi_queue_fifo_reader_in_stream_if import multi_queue_fifo_reader_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module multi_queue_fifo_reader import multi_queue_fifo_reader_pkg::*;
 (
    input wire clk,
    input wire rst,
    multi_queue_fifo_reader_in_stream_if.slave in[2],
    multi_queue_fifo_reader_out_stream_if.master out[2]
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueFifoReader
    \arq.MultiQueueFifoReader  multi_queue_fifo_reader_internal (
        .clk,
        .rst,
        .input__0__payload(in[0].p),
        .input__0__valid(in[0].valid),
        .input__0__ready(in[0].ready),
        .input__1__payload(in[1].p),
        .input__1__valid(in[1].valid),
        .input__1__ready(in[1].ready),
        .output__0__payload(out[0].p),
        .output__0__valid(out[0].valid),
        .output__0__ready(out[0].ready),
        .output__1__payload(out[1].p),
        .output__1__valid(out[1].valid),
        .output__1__ready(out[1].ready)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:892" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueFifoReader (input__0__valid, input__1__payload, input__1__valid, output__0__ready, output__1__ready, clk, rst, input__0__ready, input__1__ready, output__0__payload, output__0__valid, output__1__payload, output__1__valid, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  reg \$17 ;
  reg \$18 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:264" *)
  wire grant;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  wire input__0__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  wire input__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:262" *)
  wire next;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__0__payload;
  wire output__0__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__1__payload;
  wire output__1__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:900" *)
  reg ready_outstanding_0 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:900" *)
  reg ready_outstanding_1 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:261" *)
  wire [1:0] requests;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  assign next = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:895" *) requests;
  assign \$1  = output__0__ready | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:903" *) ready_outstanding_0;
  assign \$2  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:904" *) requests;
  assign \$3  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:904" *) grant;
  assign input__0__ready = \$2  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:904" *) \$3 ;
  assign \$4  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:905" *) ready_outstanding_0;
  assign output__0__valid = input__0__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:905" *) \$4 ;
  assign \$5  = output__1__ready | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:903" *) ready_outstanding_1;
  assign \$6  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:904" *) requests;
  assign input__1__ready = \$6  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:904" *) \$7 ;
  assign \$8  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:905" *) ready_outstanding_1;
  assign output__1__valid = input__1__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:905" *) \$8 ;
  assign \$9  = output__0__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:909" *) output__0__ready;
  assign \$10  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:909" *) input__0__ready;
  assign \$11  = \$9  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:909" *) \$10 ;
  assign \$12  = ready_outstanding_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:912" *) input__0__ready;
  assign \$13  = output__1__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:909" *) output__1__ready;
  assign \$14  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:909" *) input__1__ready;
  assign \$15  = \$13  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:909" *) \$14 ;
  assign \$16  = ready_outstanding_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:912" *) input__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:900" *)
  always @(posedge clk)
    ready_outstanding_0 <= \$17 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:900" *)
  always @(posedge clk)
    ready_outstanding_1 <= \$18 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:894" *)
  \arq.MultiQueueFifoReader.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$17  = ready_outstanding_0;
    if (\$11 ) begin
      \$17  = 1'h1;
    end
    if (\$12 ) begin
      \$17  = 1'h0;
    end
    if (rst) begin
      \$17  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$18  = ready_outstanding_1;
    if (\$15 ) begin
      \$18  = 1'h1;
    end
    if (\$16 ) begin
      \$18  = 1'h0;
    end
    if (rst) begin
      \$18  = 1'h0;
    end
  end
  assign output__0__payload = input__0__payload;
  assign output__1__payload = input__1__payload;
  assign requests[1] = \$5 ;
  assign requests[0] = \$1 ;
  assign \$7  = grant;
endmodule

(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:268" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueFifoReader.arbiter (rst, next, requests, grant, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$2  = 0;
  reg \$1 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:264" *)
  output grant;
  reg grant;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:263" *)
  reg grant_store = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:262" *)
  input next;
  wire next;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:261" *)
  input [1:0] requests;
  wire [1:0] requests;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:263" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    grant = 1'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      1'h0:
        begin
          if (requests[0]) begin
            grant = 1'h0;
          end
          if (requests[1]) begin
            grant = 1'h1;
          end
        end
      1'h1:
        begin
          if (requests[1]) begin
            grant = 1'h1;
          end
          if (requests[0]) begin
            grant = 1'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 1'h0;
    end
  end
endmodule


package cardinal_port_pkg;
typedef enum logic [2: 0] {
    LOCAL = 0,
    NORTH = 1,
    SOUTH = 2,
    EAST = 3,
    WEST = 4
} cardinal_port;
endpackage

package flit_tag_pkg;
typedef enum logic [2: 0] {
    START = 0,
    TAIL = 1,
    PAYLOAD = 2,
    START_AND_END = 3,
    ARQ_ACK = 4
} flit_tag;
endpackage

package router_crossbar_pkg;
import cardinal_port_pkg::cardinal_port;
import flit_tag_pkg::flit_tag;
export cardinal_port_pkg::cardinal_port;
export flit_tag_pkg::flit_tag;
typedef struct packed {
    logic vc_id;
    cardinal_port port;
} port;

typedef logic [5: 0][1:0] flit_arqack_credit;

typedef struct packed {
    logic [57: 0] payload;
    logic is_nack;
    logic seq_is_valid;
    flit_arqack_credit credit;
} flit_arqack;

typedef struct packed {
    logic [5: 0] y;
    logic [5: 0] x;
} coordinate;

typedef struct packed {
    coordinate target;
    logic is_flow;
} routing_target;

typedef struct packed {
    logic [58: 0] payload;
    routing_target target;
} flit_start_and_end;

typedef struct packed {
    logic [71: 0] payload;
} flit_payload;

typedef struct packed {
    logic [71: 0] payload;
} flit_tail;

typedef struct packed {
    logic [58: 0] payload;
    routing_target target;
} flit_start;

typedef union packed {
    flit_arqack arq_ack;
    flit_start_and_end start_and_end;
    flit_payload payload;
    flit_tail tail;
    flit_start start;
} flit_data;

typedef struct packed {
    flit_data data;
    flit_tag tag;
} flit;

typedef struct packed {
    port target;
    logic last;
    flit flit;
} routed_flit;

typedef struct packed {
    logic vc;
    flit flit;
} flit_with_vc;
endpackage

interface routed_flit_stream_if import router_crossbar_pkg::*;;
    routed_flit payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface router_crossbar_credit_stream_if import router_crossbar_pkg::*;;
    logic [5: 0] payload[2];
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface flit_with_vc_stream_if import router_crossbar_pkg::*;;
    flit_with_vc payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface flit_stream_if import router_crossbar_pkg::*;;
    flit payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module router_crossbar import router_crossbar_pkg::*;
 (
    input wire clk,
    input wire rst,
    routed_flit_stream_if.slave inputs[10],
    router_crossbar_credit_stream_if.slave credit[10],
    flit_with_vc_stream_if.master cardinal_outputs[4],
    flit_stream_if.master local_outputs[2]
);
    // connect_rpc -exec amaranth-rpc yosys memory_mapped_router.RouterCrossbar
    \memory_mapped_router.RouterCrossbar  router_crossbar_internal (
        .clk,
        .rst,
        .inputs__0__payload(inputs[0].p),
        .inputs__0__valid(inputs[0].valid),
        .inputs__0__ready(inputs[0].ready),
        .inputs__1__payload(inputs[1].p),
        .inputs__1__valid(inputs[1].valid),
        .inputs__1__ready(inputs[1].ready),
        .inputs__2__payload(inputs[2].p),
        .inputs__2__valid(inputs[2].valid),
        .inputs__2__ready(inputs[2].ready),
        .inputs__3__payload(inputs[3].p),
        .inputs__3__valid(inputs[3].valid),
        .inputs__3__ready(inputs[3].ready),
        .inputs__4__payload(inputs[4].p),
        .inputs__4__valid(inputs[4].valid),
        .inputs__4__ready(inputs[4].ready),
        .inputs__5__payload(inputs[5].p),
        .inputs__5__valid(inputs[5].valid),
        .inputs__5__ready(inputs[5].ready),
        .inputs__6__payload(inputs[6].p),
        .inputs__6__valid(inputs[6].valid),
        .inputs__6__ready(inputs[6].ready),
        .inputs__7__payload(inputs[7].p),
        .inputs__7__valid(inputs[7].valid),
        .inputs__7__ready(inputs[7].ready),
        .inputs__8__payload(inputs[8].p),
        .inputs__8__valid(inputs[8].valid),
        .inputs__8__ready(inputs[8].ready),
        .inputs__9__payload(inputs[9].p),
        .inputs__9__valid(inputs[9].valid),
        .inputs__9__ready(inputs[9].ready),
        .credit__0__payload({<<6{credit[0].p}}),
        .credit__0__valid(credit[0].valid),
        .credit__1__payload({<<6{credit[1].p}}),
        .credit__1__valid(credit[1].valid),
        .credit__2__payload({<<6{credit[2].p}}),
        .credit__2__valid(credit[2].valid),
        .credit__3__payload({<<6{credit[3].p}}),
        .credit__3__valid(credit[3].valid),
        .credit__4__payload({<<6{credit[4].p}}),
        .credit__4__valid(credit[4].valid),
        .credit__5__payload({<<6{credit[5].p}}),
        .credit__5__valid(credit[5].valid),
        .credit__6__payload({<<6{credit[6].p}}),
        .credit__6__valid(credit[6].valid),
        .credit__7__payload({<<6{credit[7].p}}),
        .credit__7__valid(credit[7].valid),
        .credit__8__payload({<<6{credit[8].p}}),
        .credit__8__valid(credit[8].valid),
        .credit__9__payload({<<6{credit[9].p}}),
        .credit__9__valid(credit[9].valid),
        .cardinal_outputs__0__payload(cardinal_outputs[0].p),
        .cardinal_outputs__0__valid(cardinal_outputs[0].valid),
        .cardinal_outputs__0__ready(cardinal_outputs[0].ready),
        .cardinal_outputs__1__payload(cardinal_outputs[1].p),
        .cardinal_outputs__1__valid(cardinal_outputs[1].valid),
        .cardinal_outputs__1__ready(cardinal_outputs[1].ready),
        .cardinal_outputs__2__payload(cardinal_outputs[2].p),
        .cardinal_outputs__2__valid(cardinal_outputs[2].valid),
        .cardinal_outputs__2__ready(cardinal_outputs[2].ready),
        .cardinal_outputs__3__payload(cardinal_outputs[3].p),
        .cardinal_outputs__3__valid(cardinal_outputs[3].valid),
        .cardinal_outputs__3__ready(cardinal_outputs[3].ready),
        .local_outputs__0__payload(local_outputs[0].p),
        .local_outputs__0__valid(local_outputs[0].valid),
        .local_outputs__0__ready(local_outputs[0].ready),
        .local_outputs__1__payload(local_outputs[1].p),
        .local_outputs__1__valid(local_outputs[1].valid),
        .local_outputs__1__ready(local_outputs[1].ready)
    );

    assign credit[0].ready = 1'd1;
    assign credit[1].ready = 1'd1;
    assign credit[2].ready = 1'd1;
    assign credit[3].ready = 1'd1;
    assign credit[4].ready = 1'd1;
    assign credit[5].ready = 1'd1;
    assign credit[6].ready = 1'd1;
    assign credit[7].ready = 1'd1;
    assign credit[8].ready = 1'd1;
    assign credit[9].ready = 1'd1;
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post114, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:564" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar (inputs__0__valid, inputs__1__payload, inputs__1__valid, inputs__2__payload, inputs__2__valid, inputs__3__payload, inputs__3__valid, inputs__4__payload, inputs__4__valid, inputs__5__payload, inputs__5__valid, inputs__6__payload, inputs__6__valid, inputs__7__payload, inputs__7__valid, inputs__8__payload, inputs__8__valid, inputs__9__payload, inputs__9__valid, credit__0__payload, credit__0__valid
, credit__1__payload, credit__1__valid, credit__2__payload, credit__2__valid, credit__3__payload, credit__3__valid, credit__4__payload, credit__4__valid, credit__5__payload, credit__5__valid, credit__6__payload, credit__6__valid, credit__7__payload, credit__7__valid, credit__8__payload, credit__8__valid, credit__9__payload, credit__9__valid, cardinal_outputs__0__ready, cardinal_outputs__1__ready, cardinal_outputs__2__ready
, cardinal_outputs__3__ready, local_outputs__0__ready, local_outputs__1__ready, clk, rst, inputs__0__ready, inputs__1__ready, inputs__2__ready, inputs__3__ready, inputs__4__ready, inputs__5__ready, inputs__6__ready, inputs__7__ready, inputs__8__ready, inputs__9__ready, cardinal_outputs__0__payload, cardinal_outputs__0__valid, cardinal_outputs__1__payload, cardinal_outputs__1__valid, cardinal_outputs__2__payload, cardinal_outputs__2__valid
, cardinal_outputs__3__payload, cardinal_outputs__3__valid, local_outputs__0__payload, local_outputs__0__valid, local_outputs__1__payload, local_outputs__1__valid, inputs__0__payload);
  wire [1:0] \$1 ;
  wire [1:0] \$10 ;
  wire [2:0] \$11 ;
  wire [3:0] \$12 ;
  wire [4:0] \$13 ;
  wire [5:0] \$14 ;
  wire [1:0] \$15 ;
  wire [2:0] \$16 ;
  wire [3:0] \$17 ;
  wire [4:0] \$18 ;
  wire [5:0] \$19 ;
  wire [2:0] \$2 ;
  wire [1:0] \$20 ;
  wire [2:0] \$21 ;
  wire [3:0] \$22 ;
  wire [4:0] \$23 ;
  wire [5:0] \$24 ;
  wire [3:0] \$3 ;
  wire [4:0] \$4 ;
  wire [1:0] \$5 ;
  wire [2:0] \$6 ;
  wire [3:0] \$7 ;
  wire [4:0] \$8 ;
  wire [5:0] \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] cardinal_outputs__0__payload;
  wire [75:0] cardinal_outputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \cardinal_outputs__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input cardinal_outputs__0__ready;
  wire cardinal_outputs__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output cardinal_outputs__0__valid;
  wire cardinal_outputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] cardinal_outputs__1__payload;
  wire [75:0] cardinal_outputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \cardinal_outputs__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input cardinal_outputs__1__ready;
  wire cardinal_outputs__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output cardinal_outputs__1__valid;
  wire cardinal_outputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] cardinal_outputs__2__payload;
  wire [75:0] cardinal_outputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \cardinal_outputs__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input cardinal_outputs__2__ready;
  wire cardinal_outputs__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output cardinal_outputs__2__valid;
  wire cardinal_outputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] cardinal_outputs__3__payload;
  wire [75:0] cardinal_outputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \cardinal_outputs__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input cardinal_outputs__3__ready;
  wire cardinal_outputs__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output cardinal_outputs__3__valid;
  wire cardinal_outputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__0__payload;
  wire [11:0] credit__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] \credit__0__payload$70 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__0__payload$70[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__0__payload$70[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__0__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__0__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__0__valid;
  wire credit__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \credit__0__valid$71 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__1__payload;
  wire [11:0] credit__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] \credit__1__payload$72 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__1__payload$72[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__1__payload$72[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__1__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__1__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__1__valid;
  wire credit__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \credit__1__valid$73 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__2__payload;
  wire [11:0] credit__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] \credit__2__payload$74 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__2__payload$74[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__2__payload$74[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__2__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__2__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__2__valid;
  wire credit__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \credit__2__valid$75 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__3__payload;
  wire [11:0] credit__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] \credit__3__payload$76 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__3__payload$76[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__3__payload$76[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__3__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__3__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__3__valid;
  wire credit__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \credit__3__valid$77 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__4__payload;
  wire [11:0] credit__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__4__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__4__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__4__valid;
  wire credit__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__5__payload;
  wire [11:0] credit__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__5__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__5__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__5__valid;
  wire credit__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__6__payload;
  wire [11:0] credit__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__6__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__6__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__6__valid;
  wire credit__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__7__payload;
  wire [11:0] credit__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__7__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__7__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__7__valid;
  wire credit__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__8__payload;
  wire [11:0] credit__8__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__8__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__8__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__8__valid;
  wire credit__8__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit__9__payload;
  wire [11:0] credit__9__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__9__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__9__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit__9__valid;
  wire credit__9__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [79:0] east__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \east__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [3:0] \east__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [2:0] \east__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \east__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire east__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire east__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__0__payload$128 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$128.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload$128.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload$128.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$128.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__0__payload$162 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$162.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload$162.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload$162.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$162.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__0__payload$196 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$196.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload$196.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload$196.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$196.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__0__payload$230 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$230.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload$230.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload$230.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload$230.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$130 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$164 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$198 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$232 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$125 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$159 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$193 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$227 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__1__payload$142 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$142.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload$142.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload$142.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$142.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__1__payload$176 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$176.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload$176.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload$176.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$176.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__1__payload$210 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$210.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload$210.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload$210.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$210.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \input__1__payload$244 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$244.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload$244.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload$244.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload$244.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$144 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$178 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$212 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$246 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$139 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$173 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$207 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$241 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$119 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$133 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$153 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$167 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$187 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$201 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$221 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$235 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__ready$99 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$118 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$132 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$152 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$166 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$186 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$200 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$220 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$234 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__valid$98 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  wire [3:0] input_ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  wire [3:0] \input_ready$339 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  wire [3:0] \input_ready$340 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  wire [3:0] \input_ready$341 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  wire [3:0] \input_ready$342 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  wire [3:0] \input_ready$343 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__0__payload;
  wire [79:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__0__payload$248 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$248.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload$248.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload$248.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$248.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__0__payload$263 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$263.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload$263.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload$263.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$263.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__0__payload$278 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$278.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload$278.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload$278.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$278.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__0__payload$293 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$293.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload$293.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload$293.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$293.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__0__payload$308 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$308.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload$308.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload$308.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$308.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__0__payload$323 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$323.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload$323.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload$323.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$323.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__0__payload$88 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$88.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload$88.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload$88.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload$88.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__0__ready;
  wire inputs__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__0__ready$249 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__0__ready$264 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__0__ready$279 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__0__ready$294 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__0__ready$309 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__0__ready$324 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__0__ready$90 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__0__valid$250 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__0__valid$265 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__0__valid$280 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__0__valid$295 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__0__valid$310 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__0__valid$325 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__0__valid$86 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__1__payload;
  wire [79:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__1__payload$102 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$102.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload$102.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload$102.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$102.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__1__payload$251 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$251.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload$251.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload$251.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$251.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__1__payload$266 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$266.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload$266.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload$266.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$266.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__1__payload$281 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$281.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload$281.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload$281.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$281.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__1__payload$296 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$296.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload$296.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload$296.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$296.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__1__payload$311 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$311.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload$311.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload$311.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$311.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__1__payload$326 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$326.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload$326.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload$326.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload$326.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__1__ready;
  wire inputs__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__1__ready$104 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__1__ready$252 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__1__ready$267 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__1__ready$282 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__1__ready$297 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__1__ready$312 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__1__ready$327 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__1__valid$100 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__1__valid$253 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__1__valid$268 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__1__valid$283 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__1__valid$298 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__1__valid$313 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__1__valid$328 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__2__payload;
  wire [79:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__2__payload$122 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$122.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload$122.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload$122.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$122.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__2__payload$254 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$254.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload$254.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload$254.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$254.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__2__payload$269 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$269.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload$269.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload$269.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$269.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__2__payload$284 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$284.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload$284.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload$284.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$284.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__2__payload$299 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$299.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload$299.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload$299.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$299.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__2__payload$314 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$314.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload$314.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload$314.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$314.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__2__payload$329 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$329.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload$329.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload$329.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload$329.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__2__ready;
  wire inputs__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__2__ready$124 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__2__ready$255 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__2__ready$270 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__2__ready$285 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__2__ready$300 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__2__ready$315 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__2__ready$330 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__2__valid$120 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__2__valid$256 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__2__valid$271 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__2__valid$286 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__2__valid$301 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__2__valid$316 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__2__valid$331 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__3__payload;
  wire [79:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__3__payload$136 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$136.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload$136.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload$136.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$136.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__3__payload$257 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$257.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload$257.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload$257.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$257.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__3__payload$272 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$272.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload$272.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload$272.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$272.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__3__payload$287 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$287.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload$287.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload$287.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$287.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__3__payload$302 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$302.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload$302.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload$302.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$302.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__3__payload$317 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$317.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload$317.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload$317.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$317.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [79:0] \inputs__3__payload$332 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$332.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload$332.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload$332.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload$332.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__3__ready;
  wire inputs__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__3__ready$138 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__3__ready$258 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__3__ready$273 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__3__ready$288 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__3__ready$303 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__3__ready$318 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__3__ready$333 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__3__valid$134 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__3__valid$259 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__3__valid$274 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__3__valid$289 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__3__valid$304 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__3__valid$319 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__3__valid$334 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__4__payload;
  wire [79:0] inputs__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__4__payload$156 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__4__payload$156.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__4__payload$156.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__4__payload$156.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__4__payload$156.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__4__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__4__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__4__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__4__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__4__ready;
  wire inputs__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__4__ready$158 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__4__valid;
  wire inputs__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__4__valid$154 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__5__payload;
  wire [79:0] inputs__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__5__payload$170 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__5__payload$170.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__5__payload$170.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__5__payload$170.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__5__payload$170.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__5__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__5__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__5__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__5__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__5__ready;
  wire inputs__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__5__ready$172 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__5__valid;
  wire inputs__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__5__valid$168 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__6__payload;
  wire [79:0] inputs__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__6__payload$190 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__6__payload$190.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__6__payload$190.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__6__payload$190.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__6__payload$190.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__6__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__6__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__6__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__6__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__6__ready;
  wire inputs__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__6__ready$192 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__6__valid;
  wire inputs__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__6__valid$188 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__7__payload;
  wire [79:0] inputs__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__7__payload$204 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__7__payload$204.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__7__payload$204.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__7__payload$204.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__7__payload$204.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__7__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__7__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__7__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__7__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__7__ready;
  wire inputs__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__7__ready$206 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__7__valid;
  wire inputs__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__7__valid$202 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__8__payload;
  wire [79:0] inputs__8__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__8__payload$224 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__8__payload$224.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__8__payload$224.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__8__payload$224.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__8__payload$224.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__8__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__8__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__8__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__8__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__8__ready;
  wire inputs__8__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__8__ready$226 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__8__valid;
  wire inputs__8__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__8__valid$222 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__9__payload;
  wire [79:0] inputs__9__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [4:0] \inputs__9__payload$238 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__9__payload$238.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__9__payload$238.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__9__payload$238.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__9__payload$238.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__9__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__9__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__9__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__9__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__9__ready;
  wire inputs__9__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \inputs__9__ready$240 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__9__valid;
  wire inputs__9__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \inputs__9__valid$236 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [79:0] local__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \local__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [3:0] \local__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [2:0] \local__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \local__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire local__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire local__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  output [74:0] local_outputs__0__payload;
  wire [74:0] local_outputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input local_outputs__0__ready;
  wire local_outputs__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output local_outputs__0__valid;
  wire local_outputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  output [74:0] local_outputs__1__payload;
  wire [74:0] local_outputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input local_outputs__1__ready;
  wire local_outputs__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output local_outputs__1__valid;
  wire local_outputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [79:0] north__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \north__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [3:0] \north__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [2:0] \north__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \north__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire north__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire north__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$103 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$123 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$137 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$157 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$171 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$191 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$205 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$225 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__0__ready$239 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$101 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$121 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$135 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$155 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$169 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$189 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$203 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$223 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$237 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$111 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$131 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$145 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$165 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$179 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$199 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$213 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$233 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__1__ready$247 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$107 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$127 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$141 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$161 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$175 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$195 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$209 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$229 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$243 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [80:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [80:0] \output__payload$115 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload$115.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$115.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload$115.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload$115.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$115.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$115.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [80:0] \output__payload$149 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload$149.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$149.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload$149.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload$149.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$149.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$149.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [80:0] \output__payload$183 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload$183.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$183.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload$183.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload$183.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$183.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$183.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [80:0] \output__payload$217 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload$217.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$217.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload$217.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload$217.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$217.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$217.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire [75:0] \output__payload$260 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload$260.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire [75:0] \output__payload$275 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload$275.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire [75:0] \output__payload$290 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload$290.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire [75:0] \output__payload$305 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload$305.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire [75:0] \output__payload$321 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload$321.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire [75:0] \output__payload$336 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload$336.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$116 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$150 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$184 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$218 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$261 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$276 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$291 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$306 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$322 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$337 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$113 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$147 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$181 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$215 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$262 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$277 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$292 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$307 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$320 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$335 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__8__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__8__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire outputs__9__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire outputs__9__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [79:0] south__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \south__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [3:0] \south__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [2:0] \south__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \south__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire south__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire south__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [79:0] west__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \west__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [3:0] \west__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire [2:0] \west__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:576" *)
  wire \west__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire west__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire west__valid;
  assign input__0__valid = outputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) output__1__valid;
  assign outputs__0__ready = input__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) output__1__valid;
  assign output__1__ready = input__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__0__valid;
  assign input__1__valid = outputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$107 ;
  assign outputs__1__ready = input__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$107 ;
  assign \output__1__ready$111  = input__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__1__valid;
  assign \input__0__valid$125  = outputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$127 ;
  assign outputs__2__ready = \input__0__ready$130  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$127 ;
  assign \output__1__ready$131  = \input__0__ready$130  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__2__valid;
  assign \input__1__valid$139  = outputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$141 ;
  assign outputs__3__ready = \input__1__ready$144  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$141 ;
  assign \output__1__ready$145  = \input__1__ready$144  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__3__valid;
  assign \input__0__valid$159  = outputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$161 ;
  assign outputs__4__ready = \input__0__ready$164  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$161 ;
  assign \output__1__ready$165  = \input__0__ready$164  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__4__valid;
  assign \input__1__valid$173  = outputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$175 ;
  assign outputs__5__ready = \input__1__ready$178  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$175 ;
  assign \output__1__ready$179  = \input__1__ready$178  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__5__valid;
  assign \input__0__valid$193  = outputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$195 ;
  assign outputs__6__ready = \input__0__ready$198  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$195 ;
  assign \output__1__ready$199  = \input__0__ready$198  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__6__valid;
  assign \input__1__valid$207  = outputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$209 ;
  assign outputs__7__ready = \input__1__ready$212  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$209 ;
  assign \output__1__ready$213  = \input__1__ready$212  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__7__valid;
  assign \input__0__valid$227  = outputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$229 ;
  assign outputs__8__ready = \input__0__ready$232  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$229 ;
  assign \output__1__ready$233  = \input__0__ready$232  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__8__valid;
  assign \input__1__valid$241  = outputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:605" *) \output__1__valid$243 ;
  assign outputs__9__ready = \input__1__ready$246  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:608" *) \output__1__valid$243 ;
  assign \output__1__ready$247  = \input__1__ready$246  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:609" *) outputs__9__valid;
  assign \$1  = 1'h0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) input_ready[0];
  assign \$2  = \$1  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$339 [0];
  assign \$3  = \$2  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$340 [0];
  assign \$4  = \$3  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$341 [0];
  assign \$5  = 1'h0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$339 [1];
  assign \$6  = \$5  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$340 [1];
  assign \$7  = \$6  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$341 [1];
  assign \$8  = \$7  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$342 [0];
  assign \$9  = \$8  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$343 [0];
  assign \$10  = 1'h0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) input_ready[1];
  assign \$11  = \$10  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$340 [2];
  assign \$12  = \$11  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$341 [2];
  assign \$13  = \$12  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$342 [1];
  assign \$14  = \$13  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$343 [1];
  assign \$15  = 1'h0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) input_ready[2];
  assign \$16  = \$15  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$339 [2];
  assign \$17  = \$16  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$341 [3];
  assign \$18  = \$17  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$342 [2];
  assign \$19  = \$18  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$343 [2];
  assign \$20  = 1'h0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) input_ready[3];
  assign \$21  = \$20  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$339 [3];
  assign \$22  = \$21  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$340 [3];
  assign \$23  = \$22  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$342 [3];
  assign \$24  = \$23  + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:628" *) \input_ready$343 [3];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:574" *)
  \memory_mapped_router.RouterCrossbar.crossbar_east_arb  crossbar_east_arb (
    .clk(clk),
    .input__0__payload(inputs__6__payload),
    .input__0__ready(\input__0__ready$198 ),
    .input__0__valid(\input__0__valid$193 ),
    .input__1__payload(inputs__7__payload),
    .input__1__ready(\input__1__ready$212 ),
    .input__1__valid(\input__1__valid$207 ),
    .output__payload(\output__payload$183 ),
    .output__ready(\$19 [0]),
    .output__valid(east__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_east_vc_0_tee  crossbar_east_vc_0_tee (
    .clk(clk),
    .input__ready(inputs__6__ready),
    .input__valid(inputs__6__valid),
    .output__0__ready(\output__0__ready$191 ),
    .output__0__valid(\inputs__6__valid$188 ),
    .output__1__ready(\output__1__ready$199 ),
    .output__1__valid(\output__1__valid$195 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_east_vc_1_tee  crossbar_east_vc_1_tee (
    .clk(clk),
    .input__ready(inputs__7__ready),
    .input__valid(inputs__7__valid),
    .output__0__ready(\output__0__ready$205 ),
    .output__0__valid(\inputs__7__valid$202 ),
    .output__1__ready(\output__1__ready$213 ),
    .output__1__valid(\output__1__valid$209 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:574" *)
  \memory_mapped_router.RouterCrossbar.crossbar_local_arb  crossbar_local_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload),
    .input__0__ready(input__0__ready),
    .input__0__valid(input__0__valid),
    .input__1__payload(inputs__1__payload),
    .input__1__ready(input__1__ready),
    .input__1__valid(input__1__valid),
    .output__payload(output__payload),
    .output__ready(\$4 [0]),
    .output__valid(local__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_local_vc_0_tee  crossbar_local_vc_0_tee (
    .clk(clk),
    .input__ready(inputs__0__ready),
    .input__valid(inputs__0__valid),
    .output__0__ready(output__0__ready),
    .output__0__valid(\inputs__0__valid$86 ),
    .output__1__ready(output__1__ready),
    .output__1__valid(output__1__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_local_vc_1_tee  crossbar_local_vc_1_tee (
    .clk(clk),
    .input__ready(inputs__1__ready),
    .input__valid(inputs__1__valid),
    .output__0__ready(\output__0__ready$103 ),
    .output__0__valid(\inputs__1__valid$100 ),
    .output__1__ready(\output__1__ready$111 ),
    .output__1__valid(\output__1__valid$107 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:574" *)
  \memory_mapped_router.RouterCrossbar.crossbar_north_arb  crossbar_north_arb (
    .clk(clk),
    .input__0__payload(inputs__2__payload),
    .input__0__ready(\input__0__ready$130 ),
    .input__0__valid(\input__0__valid$125 ),
    .input__1__payload(inputs__3__payload),
    .input__1__ready(\input__1__ready$144 ),
    .input__1__valid(\input__1__valid$139 ),
    .output__payload(\output__payload$115 ),
    .output__ready(\$9 [0]),
    .output__valid(north__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_north_vc_0_tee  crossbar_north_vc_0_tee (
    .clk(clk),
    .input__ready(inputs__2__ready),
    .input__valid(inputs__2__valid),
    .output__0__ready(\output__0__ready$123 ),
    .output__0__valid(\inputs__2__valid$120 ),
    .output__1__ready(\output__1__ready$131 ),
    .output__1__valid(\output__1__valid$127 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_north_vc_1_tee  crossbar_north_vc_1_tee (
    .clk(clk),
    .input__ready(inputs__3__ready),
    .input__valid(inputs__3__valid),
    .output__0__ready(\output__0__ready$137 ),
    .output__0__valid(\inputs__3__valid$134 ),
    .output__1__ready(\output__1__ready$145 ),
    .output__1__valid(\output__1__valid$141 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:617" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_east  crossbar_output_east (
    .clk(clk),
    .input_ready(\input_ready$340 ),
    .inputs__0__payload(output__payload[79:0]),
    .inputs__0__valid(local__valid),
    .inputs__1__payload(\output__payload$115 [79:0]),
    .inputs__1__valid(north__valid),
    .inputs__2__payload(\output__payload$149 [79:0]),
    .inputs__2__valid(south__valid),
    .inputs__3__payload(\output__payload$217 [79:0]),
    .inputs__3__valid(west__valid),
    .output__payload(cardinal_outputs__2__payload),
    .output__ready(cardinal_outputs__2__ready),
    .output__valid(cardinal_outputs__2__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:617" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_0  crossbar_output_local_vc_0 (
    .clk(clk),
    .input_ready(\input_ready$342 ),
    .inputs__0__payload(\output__payload$115 [79:0]),
    .inputs__0__valid(north__valid),
    .inputs__1__payload(\output__payload$149 [79:0]),
    .inputs__1__valid(south__valid),
    .inputs__2__payload(\output__payload$183 [79:0]),
    .inputs__2__valid(east__valid),
    .inputs__3__payload(\output__payload$217 [79:0]),
    .inputs__3__valid(west__valid),
    .output__payload(\output__payload$321 ),
    .output__ready(local_outputs__0__ready),
    .output__valid(local_outputs__0__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:617" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_1  crossbar_output_local_vc_1 (
    .clk(clk),
    .input_ready(\input_ready$343 ),
    .inputs__0__payload(\output__payload$115 [79:0]),
    .inputs__0__valid(north__valid),
    .inputs__1__payload(\output__payload$149 [79:0]),
    .inputs__1__valid(south__valid),
    .inputs__2__payload(\output__payload$183 [79:0]),
    .inputs__2__valid(east__valid),
    .inputs__3__payload(\output__payload$217 [79:0]),
    .inputs__3__valid(west__valid),
    .output__payload(\output__payload$336 ),
    .output__ready(local_outputs__1__ready),
    .output__valid(local_outputs__1__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:617" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_north  crossbar_output_north (
    .clk(clk),
    .input_ready(input_ready),
    .inputs__0__payload(output__payload[79:0]),
    .inputs__0__valid(local__valid),
    .inputs__1__payload(\output__payload$149 [79:0]),
    .inputs__1__valid(south__valid),
    .inputs__2__payload(\output__payload$183 [79:0]),
    .inputs__2__valid(east__valid),
    .inputs__3__payload(\output__payload$217 [79:0]),
    .inputs__3__valid(west__valid),
    .output__payload(cardinal_outputs__0__payload),
    .output__ready(cardinal_outputs__0__ready),
    .output__valid(cardinal_outputs__0__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:617" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_south  crossbar_output_south (
    .clk(clk),
    .input_ready(\input_ready$339 ),
    .inputs__0__payload(output__payload[79:0]),
    .inputs__0__valid(local__valid),
    .inputs__1__payload(\output__payload$115 [79:0]),
    .inputs__1__valid(north__valid),
    .inputs__2__payload(\output__payload$183 [79:0]),
    .inputs__2__valid(east__valid),
    .inputs__3__payload(\output__payload$217 [79:0]),
    .inputs__3__valid(west__valid),
    .output__payload(cardinal_outputs__1__payload),
    .output__ready(cardinal_outputs__1__ready),
    .output__valid(cardinal_outputs__1__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:617" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_west  crossbar_output_west (
    .clk(clk),
    .input_ready(\input_ready$341 ),
    .inputs__0__payload(output__payload[79:0]),
    .inputs__0__valid(local__valid),
    .inputs__1__payload(\output__payload$115 [79:0]),
    .inputs__1__valid(north__valid),
    .inputs__2__payload(\output__payload$149 [79:0]),
    .inputs__2__valid(south__valid),
    .inputs__3__payload(\output__payload$183 [79:0]),
    .inputs__3__valid(east__valid),
    .output__payload(cardinal_outputs__3__payload),
    .output__ready(cardinal_outputs__3__ready),
    .output__valid(cardinal_outputs__3__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:574" *)
  \memory_mapped_router.RouterCrossbar.crossbar_south_arb  crossbar_south_arb (
    .clk(clk),
    .input__0__payload(inputs__4__payload),
    .input__0__ready(\input__0__ready$164 ),
    .input__0__valid(\input__0__valid$159 ),
    .input__1__payload(inputs__5__payload),
    .input__1__ready(\input__1__ready$178 ),
    .input__1__valid(\input__1__valid$173 ),
    .output__payload(\output__payload$149 ),
    .output__ready(\$14 [0]),
    .output__valid(south__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_south_vc_0_tee  crossbar_south_vc_0_tee (
    .clk(clk),
    .input__ready(inputs__4__ready),
    .input__valid(inputs__4__valid),
    .output__0__ready(\output__0__ready$157 ),
    .output__0__valid(\inputs__4__valid$154 ),
    .output__1__ready(\output__1__ready$165 ),
    .output__1__valid(\output__1__valid$161 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_south_vc_1_tee  crossbar_south_vc_1_tee (
    .clk(clk),
    .input__ready(inputs__5__ready),
    .input__valid(inputs__5__valid),
    .output__0__ready(\output__0__ready$171 ),
    .output__0__valid(\inputs__5__valid$168 ),
    .output__1__ready(\output__1__ready$179 ),
    .output__1__valid(\output__1__valid$175 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:574" *)
  \memory_mapped_router.RouterCrossbar.crossbar_west_arb  crossbar_west_arb (
    .clk(clk),
    .input__0__payload(inputs__8__payload),
    .input__0__ready(\input__0__ready$232 ),
    .input__0__valid(\input__0__valid$227 ),
    .input__1__payload(inputs__9__payload),
    .input__1__ready(\input__1__ready$246 ),
    .input__1__valid(\input__1__valid$241 ),
    .output__payload(\output__payload$217 ),
    .output__ready(\$24 [0]),
    .output__valid(west__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_west_vc_0_tee  crossbar_west_vc_0_tee (
    .clk(clk),
    .input__ready(inputs__8__ready),
    .input__valid(inputs__8__valid),
    .output__0__ready(\output__0__ready$225 ),
    .output__0__valid(\inputs__8__valid$222 ),
    .output__1__ready(\output__1__ready$233 ),
    .output__1__valid(\output__1__valid$229 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:591" *)
  \memory_mapped_router.RouterCrossbar.crossbar_west_vc_1_tee  crossbar_west_vc_1_tee (
    .clk(clk),
    .input__ready(inputs__9__ready),
    .input__valid(inputs__9__valid),
    .output__0__ready(\output__0__ready$239 ),
    .output__0__valid(\inputs__9__valid$236 ),
    .output__1__ready(\output__1__ready$247 ),
    .output__1__valid(\output__1__valid$243 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:566" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator  vc_allocator (
    .clk(clk),
    .credit_in__payload(credit__0__payload),
    .\credit_in__payload$354 (credit__1__payload),
    .\credit_in__payload$368 (credit__2__payload),
    .\credit_in__payload$382 (credit__3__payload),
    .credit_in__valid(credit__0__valid),
    .\credit_in__valid$356 (credit__1__valid),
    .\credit_in__valid$370 (credit__2__valid),
    .\credit_in__valid$384 (credit__3__valid),
    .inputs__0__payload(\inputs__0__payload$88 ),
    .inputs__0__ready(output__0__ready),
    .inputs__0__valid(\inputs__0__valid$86 ),
    .inputs__1__payload(\inputs__1__payload$102 ),
    .inputs__1__ready(\output__0__ready$103 ),
    .inputs__1__valid(\inputs__1__valid$100 ),
    .inputs__2__payload(\inputs__2__payload$122 ),
    .inputs__2__ready(\output__0__ready$123 ),
    .inputs__2__valid(\inputs__2__valid$120 ),
    .inputs__3__payload(\inputs__3__payload$136 ),
    .inputs__3__ready(\output__0__ready$137 ),
    .inputs__3__valid(\inputs__3__valid$134 ),
    .inputs__4__payload(\inputs__4__payload$156 ),
    .inputs__4__ready(\output__0__ready$157 ),
    .inputs__4__valid(\inputs__4__valid$154 ),
    .inputs__5__payload(\inputs__5__payload$170 ),
    .inputs__5__ready(\output__0__ready$171 ),
    .inputs__5__valid(\inputs__5__valid$168 ),
    .inputs__6__payload(\inputs__6__payload$190 ),
    .inputs__6__ready(\output__0__ready$191 ),
    .inputs__6__valid(\inputs__6__valid$188 ),
    .inputs__7__payload(\inputs__7__payload$204 ),
    .inputs__7__ready(\output__0__ready$205 ),
    .inputs__7__valid(\inputs__7__valid$202 ),
    .inputs__8__payload(\inputs__8__payload$224 ),
    .inputs__8__ready(\output__0__ready$225 ),
    .inputs__8__valid(\inputs__8__valid$222 ),
    .inputs__9__payload(\inputs__9__payload$238 ),
    .inputs__9__ready(\output__0__ready$239 ),
    .inputs__9__valid(\inputs__9__valid$236 ),
    .outputs__0__ready(outputs__0__ready),
    .outputs__0__valid(outputs__0__valid),
    .outputs__1__ready(outputs__1__ready),
    .outputs__1__valid(outputs__1__valid),
    .outputs__2__ready(outputs__2__ready),
    .outputs__2__valid(outputs__2__valid),
    .outputs__3__ready(outputs__3__ready),
    .outputs__3__valid(outputs__3__valid),
    .outputs__4__ready(outputs__4__ready),
    .outputs__4__valid(outputs__4__valid),
    .outputs__5__ready(outputs__5__ready),
    .outputs__5__valid(outputs__5__valid),
    .outputs__6__ready(outputs__6__ready),
    .outputs__6__valid(outputs__6__valid),
    .outputs__7__ready(outputs__7__ready),
    .outputs__7__valid(outputs__7__valid),
    .outputs__8__ready(outputs__8__ready),
    .outputs__8__valid(outputs__8__valid),
    .outputs__9__ready(outputs__9__ready),
    .outputs__9__valid(outputs__9__valid),
    .rst(rst)
  );
  assign \credit__0__payload$70  = credit__0__payload;
  assign \credit__0__valid$71  = credit__0__valid;
  assign \credit__1__payload$72  = credit__1__payload;
  assign \credit__1__valid$73  = credit__1__valid;
  assign \credit__2__payload$74  = credit__2__payload;
  assign \credit__2__valid$75  = credit__2__valid;
  assign \credit__3__payload$76  = credit__3__payload;
  assign \credit__3__valid$77  = credit__3__valid;
  assign output__valid = local__valid;
  assign local__payload = output__payload[79:0];
  assign output__ready = \$4 [0];
  assign local__ready = \$4 [0];
  assign input__valid = inputs__0__valid;
  assign input__ready = inputs__0__ready;
  assign output__0__valid = \inputs__0__valid$86 ;
  assign \inputs__0__ready$90  = output__0__ready;
  assign input__0__payload = inputs__0__payload;
  assign \input__valid$98  = inputs__1__valid;
  assign \input__ready$99  = inputs__1__ready;
  assign \output__0__valid$101  = \inputs__1__valid$100 ;
  assign \inputs__1__ready$104  = \output__0__ready$103 ;
  assign input__1__payload = inputs__1__payload;
  assign \output__valid$113  = north__valid;
  assign north__payload = \output__payload$115 [79:0];
  assign \output__ready$116  = \$9 [0];
  assign north__ready = \$9 [0];
  assign \input__valid$118  = inputs__2__valid;
  assign \input__ready$119  = inputs__2__ready;
  assign \output__0__valid$121  = \inputs__2__valid$120 ;
  assign \inputs__2__ready$124  = \output__0__ready$123 ;
  assign \input__0__payload$128  = inputs__2__payload;
  assign \input__valid$132  = inputs__3__valid;
  assign \input__ready$133  = inputs__3__ready;
  assign \output__0__valid$135  = \inputs__3__valid$134 ;
  assign \inputs__3__ready$138  = \output__0__ready$137 ;
  assign \input__1__payload$142  = inputs__3__payload;
  assign \output__valid$147  = south__valid;
  assign south__payload = \output__payload$149 [79:0];
  assign \output__ready$150  = \$14 [0];
  assign south__ready = \$14 [0];
  assign \input__valid$152  = inputs__4__valid;
  assign \input__ready$153  = inputs__4__ready;
  assign \output__0__valid$155  = \inputs__4__valid$154 ;
  assign \inputs__4__ready$158  = \output__0__ready$157 ;
  assign \input__0__payload$162  = inputs__4__payload;
  assign \input__valid$166  = inputs__5__valid;
  assign \input__ready$167  = inputs__5__ready;
  assign \output__0__valid$169  = \inputs__5__valid$168 ;
  assign \inputs__5__ready$172  = \output__0__ready$171 ;
  assign \input__1__payload$176  = inputs__5__payload;
  assign \output__valid$181  = east__valid;
  assign east__payload = \output__payload$183 [79:0];
  assign \output__ready$184  = \$19 [0];
  assign east__ready = \$19 [0];
  assign \input__valid$186  = inputs__6__valid;
  assign \input__ready$187  = inputs__6__ready;
  assign \output__0__valid$189  = \inputs__6__valid$188 ;
  assign \inputs__6__ready$192  = \output__0__ready$191 ;
  assign \input__0__payload$196  = inputs__6__payload;
  assign \input__valid$200  = inputs__7__valid;
  assign \input__ready$201  = inputs__7__ready;
  assign \output__0__valid$203  = \inputs__7__valid$202 ;
  assign \inputs__7__ready$206  = \output__0__ready$205 ;
  assign \input__1__payload$210  = inputs__7__payload;
  assign \output__valid$215  = west__valid;
  assign west__payload = \output__payload$217 [79:0];
  assign \output__ready$218  = \$24 [0];
  assign west__ready = \$24 [0];
  assign \input__valid$220  = inputs__8__valid;
  assign \input__ready$221  = inputs__8__ready;
  assign \output__0__valid$223  = \inputs__8__valid$222 ;
  assign \inputs__8__ready$226  = \output__0__ready$225 ;
  assign \input__0__payload$230  = inputs__8__payload;
  assign \input__valid$234  = inputs__9__valid;
  assign \input__ready$235  = inputs__9__ready;
  assign \output__0__valid$237  = \inputs__9__valid$236 ;
  assign \inputs__9__ready$240  = \output__0__ready$239 ;
  assign \input__1__payload$244  = inputs__9__payload;
  assign \inputs__0__payload$248  = output__payload[79:0];
  assign \inputs__0__ready$249  = 1'h0;
  assign \inputs__0__valid$250  = local__valid;
  assign \inputs__1__payload$251  = \output__payload$149 [79:0];
  assign \inputs__1__ready$252  = 1'h0;
  assign \inputs__1__valid$253  = south__valid;
  assign \inputs__2__payload$254  = \output__payload$183 [79:0];
  assign \inputs__2__ready$255  = 1'h0;
  assign \inputs__2__valid$256  = east__valid;
  assign \inputs__3__payload$257  = \output__payload$217 [79:0];
  assign \inputs__3__ready$258  = 1'h0;
  assign \inputs__3__valid$259  = west__valid;
  assign \output__payload$260  = cardinal_outputs__0__payload;
  assign \output__ready$261  = cardinal_outputs__0__ready;
  assign \output__valid$262  = cardinal_outputs__0__valid;
  assign \inputs__0__payload$263  = output__payload[79:0];
  assign \inputs__0__ready$264  = 1'h0;
  assign \inputs__0__valid$265  = local__valid;
  assign \inputs__1__payload$266  = \output__payload$115 [79:0];
  assign \inputs__1__ready$267  = 1'h0;
  assign \inputs__1__valid$268  = north__valid;
  assign \inputs__2__payload$269  = \output__payload$183 [79:0];
  assign \inputs__2__ready$270  = 1'h0;
  assign \inputs__2__valid$271  = east__valid;
  assign \inputs__3__payload$272  = \output__payload$217 [79:0];
  assign \inputs__3__ready$273  = 1'h0;
  assign \inputs__3__valid$274  = west__valid;
  assign \output__payload$275  = cardinal_outputs__1__payload;
  assign \output__ready$276  = cardinal_outputs__1__ready;
  assign \output__valid$277  = cardinal_outputs__1__valid;
  assign \inputs__0__payload$278  = output__payload[79:0];
  assign \inputs__0__ready$279  = 1'h0;
  assign \inputs__0__valid$280  = local__valid;
  assign \inputs__1__payload$281  = \output__payload$115 [79:0];
  assign \inputs__1__ready$282  = 1'h0;
  assign \inputs__1__valid$283  = north__valid;
  assign \inputs__2__payload$284  = \output__payload$149 [79:0];
  assign \inputs__2__ready$285  = 1'h0;
  assign \inputs__2__valid$286  = south__valid;
  assign \inputs__3__payload$287  = \output__payload$217 [79:0];
  assign \inputs__3__ready$288  = 1'h0;
  assign \inputs__3__valid$289  = west__valid;
  assign \output__payload$290  = cardinal_outputs__2__payload;
  assign \output__ready$291  = cardinal_outputs__2__ready;
  assign \output__valid$292  = cardinal_outputs__2__valid;
  assign \inputs__0__payload$293  = output__payload[79:0];
  assign \inputs__0__ready$294  = 1'h0;
  assign \inputs__0__valid$295  = local__valid;
  assign \inputs__1__payload$296  = \output__payload$115 [79:0];
  assign \inputs__1__ready$297  = 1'h0;
  assign \inputs__1__valid$298  = north__valid;
  assign \inputs__2__payload$299  = \output__payload$149 [79:0];
  assign \inputs__2__ready$300  = 1'h0;
  assign \inputs__2__valid$301  = south__valid;
  assign \inputs__3__payload$302  = \output__payload$183 [79:0];
  assign \inputs__3__ready$303  = 1'h0;
  assign \inputs__3__valid$304  = east__valid;
  assign \output__payload$305  = cardinal_outputs__3__payload;
  assign \output__ready$306  = cardinal_outputs__3__ready;
  assign \output__valid$307  = cardinal_outputs__3__valid;
  assign \inputs__0__payload$308  = \output__payload$115 [79:0];
  assign \inputs__0__ready$309  = 1'h0;
  assign \inputs__0__valid$310  = north__valid;
  assign \inputs__1__payload$311  = \output__payload$149 [79:0];
  assign \inputs__1__ready$312  = 1'h0;
  assign \inputs__1__valid$313  = south__valid;
  assign \inputs__2__payload$314  = \output__payload$183 [79:0];
  assign \inputs__2__ready$315  = 1'h0;
  assign \inputs__2__valid$316  = east__valid;
  assign \inputs__3__payload$317  = \output__payload$217 [79:0];
  assign \inputs__3__ready$318  = 1'h0;
  assign \inputs__3__valid$319  = west__valid;
  assign \output__valid$320  = local_outputs__0__valid;
  assign \output__ready$322  = local_outputs__0__ready;
  assign \inputs__0__payload$323  = \output__payload$115 [79:0];
  assign \inputs__0__ready$324  = 1'h0;
  assign \inputs__0__valid$325  = north__valid;
  assign \inputs__1__payload$326  = \output__payload$149 [79:0];
  assign \inputs__1__ready$327  = 1'h0;
  assign \inputs__1__valid$328  = south__valid;
  assign \inputs__2__payload$329  = \output__payload$183 [79:0];
  assign \inputs__2__ready$330  = 1'h0;
  assign \inputs__2__valid$331  = east__valid;
  assign \inputs__3__payload$332  = \output__payload$217 [79:0];
  assign \inputs__3__ready$333  = 1'h0;
  assign \inputs__3__valid$334  = west__valid;
  assign \output__valid$335  = local_outputs__1__valid;
  assign \output__ready$337  = local_outputs__1__ready;
  assign local_outputs__0__payload = \output__payload$321 [74:0];
  assign local_outputs__1__payload = \output__payload$336 [74:0];
  assign \inputs__0__payload.last  = inputs__0__payload[75];
  assign \inputs__0__payload.target  = inputs__0__payload[79:76];
  assign \inputs__0__payload.target.port  = inputs__0__payload[78:76];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \inputs__1__payload.last  = inputs__1__payload[75];
  assign \inputs__1__payload.target  = inputs__1__payload[79:76];
  assign \inputs__1__payload.target.port  = inputs__1__payload[78:76];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \inputs__2__payload.last  = inputs__2__payload[75];
  assign \inputs__2__payload.target  = inputs__2__payload[79:76];
  assign \inputs__2__payload.target.port  = inputs__2__payload[78:76];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[79];
  assign \inputs__3__payload.last  = inputs__3__payload[75];
  assign \inputs__3__payload.target  = inputs__3__payload[79:76];
  assign \inputs__3__payload.target.port  = inputs__3__payload[78:76];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[79];
  assign \inputs__4__payload.last  = inputs__4__payload[75];
  assign \inputs__4__payload.target  = inputs__4__payload[79:76];
  assign \inputs__4__payload.target.port  = inputs__4__payload[78:76];
  assign \inputs__4__payload.target.vc_id  = inputs__4__payload[79];
  assign \inputs__5__payload.last  = inputs__5__payload[75];
  assign \inputs__5__payload.target  = inputs__5__payload[79:76];
  assign \inputs__5__payload.target.port  = inputs__5__payload[78:76];
  assign \inputs__5__payload.target.vc_id  = inputs__5__payload[79];
  assign \inputs__6__payload.last  = inputs__6__payload[75];
  assign \inputs__6__payload.target  = inputs__6__payload[79:76];
  assign \inputs__6__payload.target.port  = inputs__6__payload[78:76];
  assign \inputs__6__payload.target.vc_id  = inputs__6__payload[79];
  assign \inputs__7__payload.last  = inputs__7__payload[75];
  assign \inputs__7__payload.target  = inputs__7__payload[79:76];
  assign \inputs__7__payload.target.port  = inputs__7__payload[78:76];
  assign \inputs__7__payload.target.vc_id  = inputs__7__payload[79];
  assign \inputs__8__payload.last  = inputs__8__payload[75];
  assign \inputs__8__payload.target  = inputs__8__payload[79:76];
  assign \inputs__8__payload.target.port  = inputs__8__payload[78:76];
  assign \inputs__8__payload.target.vc_id  = inputs__8__payload[79];
  assign \inputs__9__payload.last  = inputs__9__payload[75];
  assign \inputs__9__payload.target  = inputs__9__payload[79:76];
  assign \inputs__9__payload.target.port  = inputs__9__payload[78:76];
  assign \inputs__9__payload.target.vc_id  = inputs__9__payload[79];
  assign \credit__0__payload[0]  = credit__0__payload[5:0];
  assign \credit__0__payload[1]  = credit__0__payload[11:6];
  assign \credit__1__payload[0]  = credit__1__payload[5:0];
  assign \credit__1__payload[1]  = credit__1__payload[11:6];
  assign \credit__2__payload[0]  = credit__2__payload[5:0];
  assign \credit__2__payload[1]  = credit__2__payload[11:6];
  assign \credit__3__payload[0]  = credit__3__payload[5:0];
  assign \credit__3__payload[1]  = credit__3__payload[11:6];
  assign \credit__4__payload[0]  = credit__4__payload[5:0];
  assign \credit__4__payload[1]  = credit__4__payload[11:6];
  assign \credit__5__payload[0]  = credit__5__payload[5:0];
  assign \credit__5__payload[1]  = credit__5__payload[11:6];
  assign \credit__6__payload[0]  = credit__6__payload[5:0];
  assign \credit__6__payload[1]  = credit__6__payload[11:6];
  assign \credit__7__payload[0]  = credit__7__payload[5:0];
  assign \credit__7__payload[1]  = credit__7__payload[11:6];
  assign \credit__8__payload[0]  = credit__8__payload[5:0];
  assign \credit__8__payload[1]  = credit__8__payload[11:6];
  assign \credit__9__payload[0]  = credit__9__payload[5:0];
  assign \credit__9__payload[1]  = credit__9__payload[11:6];
  assign \cardinal_outputs__0__payload.vc  = cardinal_outputs__0__payload[75];
  assign \cardinal_outputs__1__payload.vc  = cardinal_outputs__1__payload[75];
  assign \cardinal_outputs__2__payload.vc  = cardinal_outputs__2__payload[75];
  assign \cardinal_outputs__3__payload.vc  = cardinal_outputs__3__payload[75];
  assign \credit__0__payload$70[0]  = credit__0__payload[5:0];
  assign \credit__0__payload$70[1]  = credit__0__payload[11:6];
  assign \credit__1__payload$72[0]  = credit__1__payload[5:0];
  assign \credit__1__payload$72[1]  = credit__1__payload[11:6];
  assign \credit__2__payload$74[0]  = credit__2__payload[5:0];
  assign \credit__2__payload$74[1]  = credit__2__payload[11:6];
  assign \credit__3__payload$76[0]  = credit__3__payload[5:0];
  assign \credit__3__payload$76[1]  = credit__3__payload[11:6];
  assign \local__payload.last  = output__payload[75];
  assign \local__payload.target  = output__payload[79:76];
  assign \local__payload.target.port  = output__payload[78:76];
  assign \local__payload.target.vc_id  = output__payload[79];
  assign \output__payload.p  = output__payload[79:0];
  assign \output__payload.p.last  = output__payload[75];
  assign \output__payload.p.target  = output__payload[79:76];
  assign \output__payload.p.target.port  = output__payload[78:76];
  assign \output__payload.p.target.vc_id  = output__payload[79];
  assign \output__payload.src  = output__payload[80];
  assign \inputs__0__payload$88.target  = \inputs__0__payload$88 [3:0];
  assign \inputs__0__payload$88.target.port  = \inputs__0__payload$88 [2:0];
  assign \inputs__0__payload$88.target.vc_id  = \inputs__0__payload$88 [3];
  assign \inputs__0__payload$88.last  = \inputs__0__payload$88 [4];
  assign \input__0__payload.last  = inputs__0__payload[75];
  assign \input__0__payload.target  = inputs__0__payload[79:76];
  assign \input__0__payload.target.port  = inputs__0__payload[78:76];
  assign \input__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \inputs__1__payload$102.target  = \inputs__1__payload$102 [3:0];
  assign \inputs__1__payload$102.target.port  = \inputs__1__payload$102 [2:0];
  assign \inputs__1__payload$102.target.vc_id  = \inputs__1__payload$102 [3];
  assign \inputs__1__payload$102.last  = \inputs__1__payload$102 [4];
  assign \input__1__payload.last  = inputs__1__payload[75];
  assign \input__1__payload.target  = inputs__1__payload[79:76];
  assign \input__1__payload.target.port  = inputs__1__payload[78:76];
  assign \input__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \north__payload.last  = \output__payload$115 [75];
  assign \north__payload.target  = \output__payload$115 [79:76];
  assign \north__payload.target.port  = \output__payload$115 [78:76];
  assign \north__payload.target.vc_id  = \output__payload$115 [79];
  assign \output__payload$115.p  = \output__payload$115 [79:0];
  assign \output__payload$115.p.last  = \output__payload$115 [75];
  assign \output__payload$115.p.target  = \output__payload$115 [79:76];
  assign \output__payload$115.p.target.port  = \output__payload$115 [78:76];
  assign \output__payload$115.p.target.vc_id  = \output__payload$115 [79];
  assign \output__payload$115.src  = \output__payload$115 [80];
  assign \inputs__2__payload$122.target  = \inputs__2__payload$122 [3:0];
  assign \inputs__2__payload$122.target.port  = \inputs__2__payload$122 [2:0];
  assign \inputs__2__payload$122.target.vc_id  = \inputs__2__payload$122 [3];
  assign \inputs__2__payload$122.last  = \inputs__2__payload$122 [4];
  assign \input__0__payload$128.last  = inputs__2__payload[75];
  assign \input__0__payload$128.target  = inputs__2__payload[79:76];
  assign \input__0__payload$128.target.port  = inputs__2__payload[78:76];
  assign \input__0__payload$128.target.vc_id  = inputs__2__payload[79];
  assign \inputs__3__payload$136.target  = \inputs__3__payload$136 [3:0];
  assign \inputs__3__payload$136.target.port  = \inputs__3__payload$136 [2:0];
  assign \inputs__3__payload$136.target.vc_id  = \inputs__3__payload$136 [3];
  assign \inputs__3__payload$136.last  = \inputs__3__payload$136 [4];
  assign \input__1__payload$142.last  = inputs__3__payload[75];
  assign \input__1__payload$142.target  = inputs__3__payload[79:76];
  assign \input__1__payload$142.target.port  = inputs__3__payload[78:76];
  assign \input__1__payload$142.target.vc_id  = inputs__3__payload[79];
  assign \south__payload.last  = \output__payload$149 [75];
  assign \south__payload.target  = \output__payload$149 [79:76];
  assign \south__payload.target.port  = \output__payload$149 [78:76];
  assign \south__payload.target.vc_id  = \output__payload$149 [79];
  assign \output__payload$149.p  = \output__payload$149 [79:0];
  assign \output__payload$149.p.last  = \output__payload$149 [75];
  assign \output__payload$149.p.target  = \output__payload$149 [79:76];
  assign \output__payload$149.p.target.port  = \output__payload$149 [78:76];
  assign \output__payload$149.p.target.vc_id  = \output__payload$149 [79];
  assign \output__payload$149.src  = \output__payload$149 [80];
  assign \inputs__4__payload$156.target  = \inputs__4__payload$156 [3:0];
  assign \inputs__4__payload$156.target.port  = \inputs__4__payload$156 [2:0];
  assign \inputs__4__payload$156.target.vc_id  = \inputs__4__payload$156 [3];
  assign \inputs__4__payload$156.last  = \inputs__4__payload$156 [4];
  assign \input__0__payload$162.last  = inputs__4__payload[75];
  assign \input__0__payload$162.target  = inputs__4__payload[79:76];
  assign \input__0__payload$162.target.port  = inputs__4__payload[78:76];
  assign \input__0__payload$162.target.vc_id  = inputs__4__payload[79];
  assign \inputs__5__payload$170.target  = \inputs__5__payload$170 [3:0];
  assign \inputs__5__payload$170.target.port  = \inputs__5__payload$170 [2:0];
  assign \inputs__5__payload$170.target.vc_id  = \inputs__5__payload$170 [3];
  assign \inputs__5__payload$170.last  = \inputs__5__payload$170 [4];
  assign \input__1__payload$176.last  = inputs__5__payload[75];
  assign \input__1__payload$176.target  = inputs__5__payload[79:76];
  assign \input__1__payload$176.target.port  = inputs__5__payload[78:76];
  assign \input__1__payload$176.target.vc_id  = inputs__5__payload[79];
  assign \east__payload.last  = \output__payload$183 [75];
  assign \east__payload.target  = \output__payload$183 [79:76];
  assign \east__payload.target.port  = \output__payload$183 [78:76];
  assign \east__payload.target.vc_id  = \output__payload$183 [79];
  assign \output__payload$183.p  = \output__payload$183 [79:0];
  assign \output__payload$183.p.last  = \output__payload$183 [75];
  assign \output__payload$183.p.target  = \output__payload$183 [79:76];
  assign \output__payload$183.p.target.port  = \output__payload$183 [78:76];
  assign \output__payload$183.p.target.vc_id  = \output__payload$183 [79];
  assign \output__payload$183.src  = \output__payload$183 [80];
  assign \inputs__6__payload$190.target  = \inputs__6__payload$190 [3:0];
  assign \inputs__6__payload$190.target.port  = \inputs__6__payload$190 [2:0];
  assign \inputs__6__payload$190.target.vc_id  = \inputs__6__payload$190 [3];
  assign \inputs__6__payload$190.last  = \inputs__6__payload$190 [4];
  assign \input__0__payload$196.last  = inputs__6__payload[75];
  assign \input__0__payload$196.target  = inputs__6__payload[79:76];
  assign \input__0__payload$196.target.port  = inputs__6__payload[78:76];
  assign \input__0__payload$196.target.vc_id  = inputs__6__payload[79];
  assign \inputs__7__payload$204.target  = \inputs__7__payload$204 [3:0];
  assign \inputs__7__payload$204.target.port  = \inputs__7__payload$204 [2:0];
  assign \inputs__7__payload$204.target.vc_id  = \inputs__7__payload$204 [3];
  assign \inputs__7__payload$204.last  = \inputs__7__payload$204 [4];
  assign \input__1__payload$210.last  = inputs__7__payload[75];
  assign \input__1__payload$210.target  = inputs__7__payload[79:76];
  assign \input__1__payload$210.target.port  = inputs__7__payload[78:76];
  assign \input__1__payload$210.target.vc_id  = inputs__7__payload[79];
  assign \west__payload.last  = \output__payload$217 [75];
  assign \west__payload.target  = \output__payload$217 [79:76];
  assign \west__payload.target.port  = \output__payload$217 [78:76];
  assign \west__payload.target.vc_id  = \output__payload$217 [79];
  assign \output__payload$217.p  = \output__payload$217 [79:0];
  assign \output__payload$217.p.last  = \output__payload$217 [75];
  assign \output__payload$217.p.target  = \output__payload$217 [79:76];
  assign \output__payload$217.p.target.port  = \output__payload$217 [78:76];
  assign \output__payload$217.p.target.vc_id  = \output__payload$217 [79];
  assign \output__payload$217.src  = \output__payload$217 [80];
  assign \inputs__8__payload$224.target  = \inputs__8__payload$224 [3:0];
  assign \inputs__8__payload$224.target.port  = \inputs__8__payload$224 [2:0];
  assign \inputs__8__payload$224.target.vc_id  = \inputs__8__payload$224 [3];
  assign \inputs__8__payload$224.last  = \inputs__8__payload$224 [4];
  assign \input__0__payload$230.last  = inputs__8__payload[75];
  assign \input__0__payload$230.target  = inputs__8__payload[79:76];
  assign \input__0__payload$230.target.port  = inputs__8__payload[78:76];
  assign \input__0__payload$230.target.vc_id  = inputs__8__payload[79];
  assign \inputs__9__payload$238.target  = \inputs__9__payload$238 [3:0];
  assign \inputs__9__payload$238.target.port  = \inputs__9__payload$238 [2:0];
  assign \inputs__9__payload$238.target.vc_id  = \inputs__9__payload$238 [3];
  assign \inputs__9__payload$238.last  = \inputs__9__payload$238 [4];
  assign \input__1__payload$244.last  = inputs__9__payload[75];
  assign \input__1__payload$244.target  = inputs__9__payload[79:76];
  assign \input__1__payload$244.target.port  = inputs__9__payload[78:76];
  assign \input__1__payload$244.target.vc_id  = inputs__9__payload[79];
  assign \inputs__0__payload$248.last  = output__payload[75];
  assign \inputs__0__payload$248.target  = output__payload[79:76];
  assign \inputs__0__payload$248.target.port  = output__payload[78:76];
  assign \inputs__0__payload$248.target.vc_id  = output__payload[79];
  assign \inputs__1__payload$251.last  = \output__payload$149 [75];
  assign \inputs__1__payload$251.target  = \output__payload$149 [79:76];
  assign \inputs__1__payload$251.target.port  = \output__payload$149 [78:76];
  assign \inputs__1__payload$251.target.vc_id  = \output__payload$149 [79];
  assign \inputs__2__payload$254.last  = \output__payload$183 [75];
  assign \inputs__2__payload$254.target  = \output__payload$183 [79:76];
  assign \inputs__2__payload$254.target.port  = \output__payload$183 [78:76];
  assign \inputs__2__payload$254.target.vc_id  = \output__payload$183 [79];
  assign \inputs__3__payload$257.last  = \output__payload$217 [75];
  assign \inputs__3__payload$257.target  = \output__payload$217 [79:76];
  assign \inputs__3__payload$257.target.port  = \output__payload$217 [78:76];
  assign \inputs__3__payload$257.target.vc_id  = \output__payload$217 [79];
  assign \output__payload$260.vc  = cardinal_outputs__0__payload[75];
  assign \inputs__0__payload$263.last  = output__payload[75];
  assign \inputs__0__payload$263.target  = output__payload[79:76];
  assign \inputs__0__payload$263.target.port  = output__payload[78:76];
  assign \inputs__0__payload$263.target.vc_id  = output__payload[79];
  assign \inputs__1__payload$266.last  = \output__payload$115 [75];
  assign \inputs__1__payload$266.target  = \output__payload$115 [79:76];
  assign \inputs__1__payload$266.target.port  = \output__payload$115 [78:76];
  assign \inputs__1__payload$266.target.vc_id  = \output__payload$115 [79];
  assign \inputs__2__payload$269.last  = \output__payload$183 [75];
  assign \inputs__2__payload$269.target  = \output__payload$183 [79:76];
  assign \inputs__2__payload$269.target.port  = \output__payload$183 [78:76];
  assign \inputs__2__payload$269.target.vc_id  = \output__payload$183 [79];
  assign \inputs__3__payload$272.last  = \output__payload$217 [75];
  assign \inputs__3__payload$272.target  = \output__payload$217 [79:76];
  assign \inputs__3__payload$272.target.port  = \output__payload$217 [78:76];
  assign \inputs__3__payload$272.target.vc_id  = \output__payload$217 [79];
  assign \output__payload$275.vc  = cardinal_outputs__1__payload[75];
  assign \inputs__0__payload$278.last  = output__payload[75];
  assign \inputs__0__payload$278.target  = output__payload[79:76];
  assign \inputs__0__payload$278.target.port  = output__payload[78:76];
  assign \inputs__0__payload$278.target.vc_id  = output__payload[79];
  assign \inputs__1__payload$281.last  = \output__payload$115 [75];
  assign \inputs__1__payload$281.target  = \output__payload$115 [79:76];
  assign \inputs__1__payload$281.target.port  = \output__payload$115 [78:76];
  assign \inputs__1__payload$281.target.vc_id  = \output__payload$115 [79];
  assign \inputs__2__payload$284.last  = \output__payload$149 [75];
  assign \inputs__2__payload$284.target  = \output__payload$149 [79:76];
  assign \inputs__2__payload$284.target.port  = \output__payload$149 [78:76];
  assign \inputs__2__payload$284.target.vc_id  = \output__payload$149 [79];
  assign \inputs__3__payload$287.last  = \output__payload$217 [75];
  assign \inputs__3__payload$287.target  = \output__payload$217 [79:76];
  assign \inputs__3__payload$287.target.port  = \output__payload$217 [78:76];
  assign \inputs__3__payload$287.target.vc_id  = \output__payload$217 [79];
  assign \output__payload$290.vc  = cardinal_outputs__2__payload[75];
  assign \inputs__0__payload$293.last  = output__payload[75];
  assign \inputs__0__payload$293.target  = output__payload[79:76];
  assign \inputs__0__payload$293.target.port  = output__payload[78:76];
  assign \inputs__0__payload$293.target.vc_id  = output__payload[79];
  assign \inputs__1__payload$296.last  = \output__payload$115 [75];
  assign \inputs__1__payload$296.target  = \output__payload$115 [79:76];
  assign \inputs__1__payload$296.target.port  = \output__payload$115 [78:76];
  assign \inputs__1__payload$296.target.vc_id  = \output__payload$115 [79];
  assign \inputs__2__payload$299.last  = \output__payload$149 [75];
  assign \inputs__2__payload$299.target  = \output__payload$149 [79:76];
  assign \inputs__2__payload$299.target.port  = \output__payload$149 [78:76];
  assign \inputs__2__payload$299.target.vc_id  = \output__payload$149 [79];
  assign \inputs__3__payload$302.last  = \output__payload$183 [75];
  assign \inputs__3__payload$302.target  = \output__payload$183 [79:76];
  assign \inputs__3__payload$302.target.port  = \output__payload$183 [78:76];
  assign \inputs__3__payload$302.target.vc_id  = \output__payload$183 [79];
  assign \output__payload$305.vc  = cardinal_outputs__3__payload[75];
  assign \inputs__0__payload$308.last  = \output__payload$115 [75];
  assign \inputs__0__payload$308.target  = \output__payload$115 [79:76];
  assign \inputs__0__payload$308.target.port  = \output__payload$115 [78:76];
  assign \inputs__0__payload$308.target.vc_id  = \output__payload$115 [79];
  assign \inputs__1__payload$311.last  = \output__payload$149 [75];
  assign \inputs__1__payload$311.target  = \output__payload$149 [79:76];
  assign \inputs__1__payload$311.target.port  = \output__payload$149 [78:76];
  assign \inputs__1__payload$311.target.vc_id  = \output__payload$149 [79];
  assign \inputs__2__payload$314.last  = \output__payload$183 [75];
  assign \inputs__2__payload$314.target  = \output__payload$183 [79:76];
  assign \inputs__2__payload$314.target.port  = \output__payload$183 [78:76];
  assign \inputs__2__payload$314.target.vc_id  = \output__payload$183 [79];
  assign \inputs__3__payload$317.last  = \output__payload$217 [75];
  assign \inputs__3__payload$317.target  = \output__payload$217 [79:76];
  assign \inputs__3__payload$317.target.port  = \output__payload$217 [78:76];
  assign \inputs__3__payload$317.target.vc_id  = \output__payload$217 [79];
  assign \output__payload$321.vc  = \output__payload$321 [75];
  assign \inputs__0__payload$323.last  = \output__payload$115 [75];
  assign \inputs__0__payload$323.target  = \output__payload$115 [79:76];
  assign \inputs__0__payload$323.target.port  = \output__payload$115 [78:76];
  assign \inputs__0__payload$323.target.vc_id  = \output__payload$115 [79];
  assign \inputs__1__payload$326.last  = \output__payload$149 [75];
  assign \inputs__1__payload$326.target  = \output__payload$149 [79:76];
  assign \inputs__1__payload$326.target.port  = \output__payload$149 [78:76];
  assign \inputs__1__payload$326.target.vc_id  = \output__payload$149 [79];
  assign \inputs__2__payload$329.last  = \output__payload$183 [75];
  assign \inputs__2__payload$329.target  = \output__payload$183 [79:76];
  assign \inputs__2__payload$329.target.port  = \output__payload$183 [78:76];
  assign \inputs__2__payload$329.target.vc_id  = \output__payload$183 [79];
  assign \inputs__3__payload$332.last  = \output__payload$217 [75];
  assign \inputs__3__payload$332.target  = \output__payload$217 [79:76];
  assign \inputs__3__payload$332.target.port  = \output__payload$217 [78:76];
  assign \inputs__3__payload$332.target.vc_id  = \output__payload$217 [79];
  assign \output__payload$336.vc  = \output__payload$336 [75];
  assign \inputs__9__payload$238 [4] = inputs__9__payload[75];
  assign \inputs__9__payload$238 [3:0] = inputs__9__payload[79:76];
  assign \inputs__8__payload$224 [4] = inputs__8__payload[75];
  assign \inputs__8__payload$224 [3:0] = inputs__8__payload[79:76];
  assign \inputs__7__payload$204 [4] = inputs__7__payload[75];
  assign \inputs__7__payload$204 [3:0] = inputs__7__payload[79:76];
  assign \inputs__6__payload$190 [4] = inputs__6__payload[75];
  assign \inputs__6__payload$190 [3:0] = inputs__6__payload[79:76];
  assign \inputs__5__payload$170 [4] = inputs__5__payload[75];
  assign \inputs__5__payload$170 [3:0] = inputs__5__payload[79:76];
  assign \inputs__4__payload$156 [4] = inputs__4__payload[75];
  assign \inputs__4__payload$156 [3:0] = inputs__4__payload[79:76];
  assign \inputs__3__payload$136 [4] = inputs__3__payload[75];
  assign \inputs__3__payload$136 [3:0] = inputs__3__payload[79:76];
  assign \inputs__2__payload$122 [4] = inputs__2__payload[75];
  assign \inputs__2__payload$122 [3:0] = inputs__2__payload[79:76];
  assign \inputs__1__payload$102 [4] = inputs__1__payload[75];
  assign \inputs__1__payload$102 [3:0] = inputs__1__payload[79:76];
  assign \inputs__0__payload$88 [4] = inputs__0__payload[75];
  assign \inputs__0__payload$88 [3:0] = inputs__0__payload[79:76];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_east_arb (input__1__payload, clk, rst, input__0__valid, input__1__valid, output__ready, output__valid, output__payload, input__0__ready, input__1__ready, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  reg \$1 ;
  reg [79:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__0__payload;
  wire [79:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__1__payload;
  wire [79:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [80:0] output__payload;
  reg [80:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_east_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$1  = input__0__valid;
      1'h1:
          \$1  = input__1__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$2  = input__0__payload;
      1'h1:
          \$2  = input__1__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    output__payload = 81'h000000000000000000000;
    if (transfer) begin
      output__payload[79:0] = \$2 ;
      output__payload[80] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        1'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        1'h0:
            /* empty */;
        1'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    granted = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[79:0];
  assign \output__payload.p.last  = output__payload[75];
  assign \output__payload.p.target  = output__payload[79:76];
  assign \output__payload.p.target.port  = output__payload[78:76];
  assign \output__payload.p.target.vc_id  = output__payload[79];
  assign \output__payload.src  = output__payload[80];
  assign \input__0__payload.last  = input__0__payload[75];
  assign \input__0__payload.target  = input__0__payload[79:76];
  assign \input__0__payload.target.port  = input__0__payload[78:76];
  assign \input__0__payload.target.vc_id  = input__0__payload[79];
  assign \input__1__payload.last  = input__1__payload[75];
  assign \input__1__payload.target  = input__1__payload[79:76];
  assign \input__1__payload.target.port  = input__1__payload[78:76];
  assign \input__1__payload.target.vc_id  = input__1__payload[79];
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_east_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$2  = 0;
  reg \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output grant;
  reg grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output grant_store;
  reg grant_store = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [1:0] requests;
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    grant = 1'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      1'h0:
        begin
          if (requests[0]) begin
            grant = 1'h0;
          end
          if (requests[1]) begin
            grant = 1'h1;
          end
        end
      1'h1:
        begin
          if (requests[1]) begin
            grant = 1'h1;
          end
          if (requests[0]) begin
            grant = 1'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 1'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_east_vc_0_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$3  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$3 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$3 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_east_vc_1_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$4  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$4 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$4 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_local_arb (input__1__payload, clk, rst, input__0__valid, input__1__valid, output__ready, output__valid, output__payload, input__0__ready, input__1__ready, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$5  = 0;
  reg \$1 ;
  reg [79:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__0__payload;
  wire [79:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__1__payload;
  wire [79:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [80:0] output__payload;
  reg [80:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_local_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$1  = input__0__valid;
      1'h1:
          \$1  = input__1__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$2  = input__0__payload;
      1'h1:
          \$2  = input__1__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    output__payload = 81'h000000000000000000000;
    if (transfer) begin
      output__payload[79:0] = \$2 ;
      output__payload[80] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        1'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        1'h0:
            /* empty */;
        1'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    granted = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$5 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[79:0];
  assign \output__payload.p.last  = output__payload[75];
  assign \output__payload.p.target  = output__payload[79:76];
  assign \output__payload.p.target.port  = output__payload[78:76];
  assign \output__payload.p.target.vc_id  = output__payload[79];
  assign \output__payload.src  = output__payload[80];
  assign \input__0__payload.last  = input__0__payload[75];
  assign \input__0__payload.target  = input__0__payload[79:76];
  assign \input__0__payload.target.port  = input__0__payload[78:76];
  assign \input__0__payload.target.vc_id  = input__0__payload[79];
  assign \input__1__payload.last  = input__1__payload[75];
  assign \input__1__payload.target  = input__1__payload[79:76];
  assign \input__1__payload.target.port  = input__1__payload[78:76];
  assign \input__1__payload.target.vc_id  = input__1__payload[79];
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_local_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$6  = 0;
  reg \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output grant;
  reg grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output grant_store;
  reg grant_store = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [1:0] requests;
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$6 ) begin end
    grant = 1'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      1'h0:
        begin
          if (requests[0]) begin
            grant = 1'h0;
          end
          if (requests[1]) begin
            grant = 1'h1;
          end
        end
      1'h1:
        begin
          if (requests[1]) begin
            grant = 1'h1;
          end
          if (requests[0]) begin
            grant = 1'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$6 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 1'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_local_vc_0_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$7  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$7 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$7 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_local_vc_1_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$8  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$8 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$8 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_north_arb (input__1__payload, clk, rst, input__0__valid, input__1__valid, output__ready, output__valid, output__payload, input__0__ready, input__1__ready, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$9  = 0;
  reg \$1 ;
  reg [79:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__0__payload;
  wire [79:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__1__payload;
  wire [79:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [80:0] output__payload;
  reg [80:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_north_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$1  = input__0__valid;
      1'h1:
          \$1  = input__1__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$2  = input__0__payload;
      1'h1:
          \$2  = input__1__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    output__payload = 81'h000000000000000000000;
    if (transfer) begin
      output__payload[79:0] = \$2 ;
      output__payload[80] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        1'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        1'h0:
            /* empty */;
        1'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    granted = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$9 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[79:0];
  assign \output__payload.p.last  = output__payload[75];
  assign \output__payload.p.target  = output__payload[79:76];
  assign \output__payload.p.target.port  = output__payload[78:76];
  assign \output__payload.p.target.vc_id  = output__payload[79];
  assign \output__payload.src  = output__payload[80];
  assign \input__0__payload.last  = input__0__payload[75];
  assign \input__0__payload.target  = input__0__payload[79:76];
  assign \input__0__payload.target.port  = input__0__payload[78:76];
  assign \input__0__payload.target.vc_id  = input__0__payload[79];
  assign \input__1__payload.last  = input__1__payload[75];
  assign \input__1__payload.target  = input__1__payload[79:76];
  assign \input__1__payload.target.port  = input__1__payload[78:76];
  assign \input__1__payload.target.vc_id  = input__1__payload[79];
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_north_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$10  = 0;
  reg \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output grant;
  reg grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output grant_store;
  reg grant_store = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [1:0] requests;
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$10 ) begin end
    grant = 1'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      1'h0:
        begin
          if (requests[0]) begin
            grant = 1'h0;
          end
          if (requests[1]) begin
            grant = 1'h1;
          end
        end
      1'h1:
        begin
          if (requests[1]) begin
            grant = 1'h1;
          end
          if (requests[0]) begin
            grant = 1'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$10 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 1'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_north_vc_0_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$11  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$11 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$11 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_north_vc_1_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$12  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$12 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$12 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:454" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_east (clk, rst, inputs__0__valid, inputs__0__payload, inputs__1__valid, inputs__1__payload, inputs__2__valid, inputs__2__payload, inputs__3__valid, inputs__3__payload, input_ready, output__valid, output__payload, output__ready);
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  output [3:0] input_ready;
  wire [3:0] input_ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__0__payload;
  wire [79:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__1__payload;
  wire [79:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__2__payload;
  wire [79:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__3__payload;
  wire [79:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] output__payload;
  wire [75:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [77:0] \output__payload$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload$24.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$24.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload$24.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$26 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  assign \$1  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$2  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hb;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$2 , \$1  };
  assign input__0__valid = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$3 ;
  assign \$4  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$5  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hb;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$5 , \$4  };
  assign input__1__valid = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$6 ;
  assign \$7  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$8  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hb;
  assign \$9  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$8 , \$7  };
  assign input__2__valid = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$9 ;
  assign \$10  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$11  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hb;
  assign \$12  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$11 , \$10  };
  assign input__3__valid = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:459" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_east.arbiter  arbiter (
    .clk(clk),
    .input__0__payload(input__0__payload),
    .input__0__ready(input__0__ready),
    .input__0__valid(input__0__valid),
    .input__1__payload(input__1__payload),
    .input__1__ready(input__1__ready),
    .input__1__valid(input__1__valid),
    .input__2__payload(input__2__payload),
    .input__2__ready(input__2__ready),
    .input__2__valid(input__2__valid),
    .input__3__payload(input__3__payload),
    .input__3__ready(input__3__ready),
    .input__3__valid(input__3__valid),
    .output__payload(\output__payload$24 ),
    .output__ready(output__ready),
    .output__valid(output__valid),
    .rst(rst)
  );
  assign \output__valid$22  = output__valid;
  assign \output__ready$26  = output__ready;
  assign output__payload = \output__payload$24 [75:0];
  assign \inputs__0__payload.last  = inputs__0__payload[75];
  assign \inputs__0__payload.target  = inputs__0__payload[79:76];
  assign \inputs__0__payload.target.port  = inputs__0__payload[78:76];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \inputs__1__payload.last  = inputs__1__payload[75];
  assign \inputs__1__payload.target  = inputs__1__payload[79:76];
  assign \inputs__1__payload.target.port  = inputs__1__payload[78:76];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \inputs__2__payload.last  = inputs__2__payload[75];
  assign \inputs__2__payload.target  = inputs__2__payload[79:76];
  assign \inputs__2__payload.target.port  = inputs__2__payload[78:76];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[79];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \inputs__3__payload.last  = inputs__3__payload[75];
  assign \inputs__3__payload.target  = inputs__3__payload[79:76];
  assign \inputs__3__payload.target.port  = inputs__3__payload[78:76];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[79];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign \output__payload.vc  = \output__payload$24 [75];
  assign \output__payload$24.p  = \output__payload$24 [75:0];
  assign \output__payload$24.p.vc  = \output__payload$24 [75];
  assign \output__payload$24.src  = \output__payload$24 [77:76];
  assign input__3__payload[75] = inputs__3__payload[79];
  assign input__3__payload[74:0] = inputs__3__payload[74:0];
  assign input__2__payload[75] = inputs__2__payload[79];
  assign input__2__payload[74:0] = inputs__2__payload[74:0];
  assign input__1__payload[75] = inputs__1__payload[79];
  assign input__1__payload[74:0] = inputs__1__payload[74:0];
  assign input_ready[3] = input__3__ready;
  assign input_ready[2] = input__2__ready;
  assign input_ready[1] = input__1__ready;
  assign input_ready[0] = input__0__ready;
  assign input__0__payload[75] = inputs__0__payload[79];
  assign input__0__payload[74:0] = inputs__0__payload[74:0];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_east.arbiter (clk, rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__0__payload, input__1__payload, input__2__payload, input__3__payload, output__valid, output__payload, input__0__ready, input__1__ready, input__2__ready, input__3__ready, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$13  = 0;
  reg \$1 ;
  reg [75:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [1:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg [1:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__0__payload;
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__1__payload;
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__2__payload;
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__3__payload;
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [77:0] output__payload;
  reg [77:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_east.arbiter.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$1  = input__0__valid;
      2'h1:
          \$1  = input__1__valid;
      2'h2:
          \$1  = input__2__valid;
      2'h3:
          \$1  = input__3__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$2  = input__0__payload;
      2'h1:
          \$2  = input__1__payload;
      2'h2:
          \$2  = input__2__payload;
      2'h3:
          \$2  = input__3__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    output__payload = 78'h00000000000000000000;
    if (transfer) begin
      output__payload[75:0] = \$2 ;
      output__payload[77:76] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            /* empty */;
        2'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    granted = 2'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$13 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[75:0];
  assign \output__payload.p.vc  = output__payload[75];
  assign \output__payload.src  = output__payload[77:76];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_east.arbiter.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$14  = 0;
  reg [1:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [1:0] grant;
  reg [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [1:0] grant_store;
  reg [1:0] grant_store = 2'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [3:0] requests;
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$14 ) begin end
    grant = 2'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      2'h0:
        begin
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
        end
      2'h1:
        begin
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
        end
      2'h2:
        begin
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
        end
      2'h3:
        begin
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$14 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 2'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:454" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_0 (clk, rst, inputs__0__valid, inputs__0__payload, inputs__1__valid, inputs__1__payload, inputs__2__valid, inputs__2__payload, inputs__3__valid, inputs__3__payload, input_ready, output__valid, output__payload, output__ready);
  wire \$1 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  output [3:0] input_ready;
  wire [3:0] input_ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__0__payload;
  wire [79:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__1__payload;
  wire [79:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__2__payload;
  wire [79:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__3__payload;
  wire [79:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] output__payload;
  wire [75:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [77:0] \output__payload$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload$24.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$24.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload$24.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$26 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  assign input__2__valid = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$3 ;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) inputs__3__payload[79:76];
  assign input__3__valid = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$4 ;
  assign \$1  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) inputs__0__payload[79:76];
  assign input__0__valid = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$1 ;
  assign \$2  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) inputs__1__payload[79:76];
  assign input__1__valid = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$2 ;
  assign \$3  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) inputs__2__payload[79:76];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:459" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_0.arbiter  arbiter (
    .clk(clk),
    .input__0__payload(input__0__payload),
    .input__0__ready(input__0__ready),
    .input__0__valid(input__0__valid),
    .input__1__payload(input__1__payload),
    .input__1__ready(input__1__ready),
    .input__1__valid(input__1__valid),
    .input__2__payload(input__2__payload),
    .input__2__ready(input__2__ready),
    .input__2__valid(input__2__valid),
    .input__3__payload(input__3__payload),
    .input__3__ready(input__3__ready),
    .input__3__valid(input__3__valid),
    .output__payload(\output__payload$24 ),
    .output__ready(output__ready),
    .output__valid(output__valid),
    .rst(rst)
  );
  assign \output__valid$22  = output__valid;
  assign \output__ready$26  = output__ready;
  assign output__payload = \output__payload$24 [75:0];
  assign \inputs__0__payload.last  = inputs__0__payload[75];
  assign \inputs__0__payload.target  = inputs__0__payload[79:76];
  assign \inputs__0__payload.target.port  = inputs__0__payload[78:76];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \inputs__1__payload.last  = inputs__1__payload[75];
  assign \inputs__1__payload.target  = inputs__1__payload[79:76];
  assign \inputs__1__payload.target.port  = inputs__1__payload[78:76];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \inputs__2__payload.last  = inputs__2__payload[75];
  assign \inputs__2__payload.target  = inputs__2__payload[79:76];
  assign \inputs__2__payload.target.port  = inputs__2__payload[78:76];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[79];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \inputs__3__payload.last  = inputs__3__payload[75];
  assign \inputs__3__payload.target  = inputs__3__payload[79:76];
  assign \inputs__3__payload.target.port  = inputs__3__payload[78:76];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[79];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign \output__payload.vc  = \output__payload$24 [75];
  assign \output__payload$24.p  = \output__payload$24 [75:0];
  assign \output__payload$24.p.vc  = \output__payload$24 [75];
  assign \output__payload$24.src  = \output__payload$24 [77:76];
  assign input__3__payload[75] = inputs__3__payload[79];
  assign input__3__payload[74:0] = inputs__3__payload[74:0];
  assign input__2__payload[75] = inputs__2__payload[79];
  assign input__2__payload[74:0] = inputs__2__payload[74:0];
  assign input__1__payload[75] = inputs__1__payload[79];
  assign input__1__payload[74:0] = inputs__1__payload[74:0];
  assign input_ready[3] = input__3__ready;
  assign input_ready[2] = input__2__ready;
  assign input_ready[1] = input__1__ready;
  assign input_ready[0] = input__0__ready;
  assign input__0__payload[75] = inputs__0__payload[79];
  assign input__0__payload[74:0] = inputs__0__payload[74:0];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_0.arbiter (clk, rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__0__payload, input__1__payload, input__2__payload, input__3__payload, output__valid, output__payload, input__0__ready, input__1__ready, input__2__ready, input__3__ready, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$15  = 0;
  reg \$1 ;
  reg [75:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [1:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg [1:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__0__payload;
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__1__payload;
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__2__payload;
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__3__payload;
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [77:0] output__payload;
  reg [77:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_0.arbiter.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$1  = input__0__valid;
      2'h1:
          \$1  = input__1__valid;
      2'h2:
          \$1  = input__2__valid;
      2'h3:
          \$1  = input__3__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$2  = input__0__payload;
      2'h1:
          \$2  = input__1__payload;
      2'h2:
          \$2  = input__2__payload;
      2'h3:
          \$2  = input__3__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    output__payload = 78'h00000000000000000000;
    if (transfer) begin
      output__payload[75:0] = \$2 ;
      output__payload[77:76] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            /* empty */;
        2'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    granted = 2'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$15 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[75:0];
  assign \output__payload.p.vc  = output__payload[75];
  assign \output__payload.src  = output__payload[77:76];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_0.arbiter.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$16  = 0;
  reg [1:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [1:0] grant;
  reg [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [1:0] grant_store;
  reg [1:0] grant_store = 2'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [3:0] requests;
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$16 ) begin end
    grant = 2'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      2'h0:
        begin
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
        end
      2'h1:
        begin
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
        end
      2'h2:
        begin
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
        end
      2'h3:
        begin
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$16 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 2'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:454" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_1 (clk, rst, inputs__0__valid, inputs__0__payload, inputs__1__valid, inputs__1__payload, inputs__2__valid, inputs__2__payload, inputs__3__valid, inputs__3__payload, input_ready, output__valid, output__payload, output__ready);
  wire \$1 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  output [3:0] input_ready;
  wire [3:0] input_ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__0__payload;
  wire [79:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__1__payload;
  wire [79:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__2__payload;
  wire [79:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__3__payload;
  wire [79:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] output__payload;
  wire [75:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [77:0] \output__payload$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload$24.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$24.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload$24.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$26 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  assign input__2__valid = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$3 ;
  assign \$4  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h8;
  assign input__3__valid = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$4 ;
  assign \$1  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h8;
  assign input__0__valid = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$1 ;
  assign \$2  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h8;
  assign input__1__valid = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$2 ;
  assign \$3  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h8;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:459" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_1.arbiter  arbiter (
    .clk(clk),
    .input__0__payload(input__0__payload),
    .input__0__ready(input__0__ready),
    .input__0__valid(input__0__valid),
    .input__1__payload(input__1__payload),
    .input__1__ready(input__1__ready),
    .input__1__valid(input__1__valid),
    .input__2__payload(input__2__payload),
    .input__2__ready(input__2__ready),
    .input__2__valid(input__2__valid),
    .input__3__payload(input__3__payload),
    .input__3__ready(input__3__ready),
    .input__3__valid(input__3__valid),
    .output__payload(\output__payload$24 ),
    .output__ready(output__ready),
    .output__valid(output__valid),
    .rst(rst)
  );
  assign \output__valid$22  = output__valid;
  assign \output__ready$26  = output__ready;
  assign output__payload = \output__payload$24 [75:0];
  assign \inputs__0__payload.last  = inputs__0__payload[75];
  assign \inputs__0__payload.target  = inputs__0__payload[79:76];
  assign \inputs__0__payload.target.port  = inputs__0__payload[78:76];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \inputs__1__payload.last  = inputs__1__payload[75];
  assign \inputs__1__payload.target  = inputs__1__payload[79:76];
  assign \inputs__1__payload.target.port  = inputs__1__payload[78:76];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \inputs__2__payload.last  = inputs__2__payload[75];
  assign \inputs__2__payload.target  = inputs__2__payload[79:76];
  assign \inputs__2__payload.target.port  = inputs__2__payload[78:76];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[79];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \inputs__3__payload.last  = inputs__3__payload[75];
  assign \inputs__3__payload.target  = inputs__3__payload[79:76];
  assign \inputs__3__payload.target.port  = inputs__3__payload[78:76];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[79];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign \output__payload.vc  = \output__payload$24 [75];
  assign \output__payload$24.p  = \output__payload$24 [75:0];
  assign \output__payload$24.p.vc  = \output__payload$24 [75];
  assign \output__payload$24.src  = \output__payload$24 [77:76];
  assign input__3__payload[75] = inputs__3__payload[79];
  assign input__3__payload[74:0] = inputs__3__payload[74:0];
  assign input__2__payload[75] = inputs__2__payload[79];
  assign input__2__payload[74:0] = inputs__2__payload[74:0];
  assign input__1__payload[75] = inputs__1__payload[79];
  assign input__1__payload[74:0] = inputs__1__payload[74:0];
  assign input_ready[3] = input__3__ready;
  assign input_ready[2] = input__2__ready;
  assign input_ready[1] = input__1__ready;
  assign input_ready[0] = input__0__ready;
  assign input__0__payload[75] = inputs__0__payload[79];
  assign input__0__payload[74:0] = inputs__0__payload[74:0];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_1.arbiter (clk, rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__0__payload, input__1__payload, input__2__payload, input__3__payload, output__valid, output__payload, input__0__ready, input__1__ready, input__2__ready, input__3__ready, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$17  = 0;
  reg \$1 ;
  reg [75:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [1:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg [1:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__0__payload;
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__1__payload;
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__2__payload;
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__3__payload;
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [77:0] output__payload;
  reg [77:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_1.arbiter.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$1  = input__0__valid;
      2'h1:
          \$1  = input__1__valid;
      2'h2:
          \$1  = input__2__valid;
      2'h3:
          \$1  = input__3__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$2  = input__0__payload;
      2'h1:
          \$2  = input__1__payload;
      2'h2:
          \$2  = input__2__payload;
      2'h3:
          \$2  = input__3__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    output__payload = 78'h00000000000000000000;
    if (transfer) begin
      output__payload[75:0] = \$2 ;
      output__payload[77:76] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            /* empty */;
        2'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    granted = 2'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$17 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[75:0];
  assign \output__payload.p.vc  = output__payload[75];
  assign \output__payload.src  = output__payload[77:76];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_local_vc_1.arbiter.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$18  = 0;
  reg [1:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [1:0] grant;
  reg [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [1:0] grant_store;
  reg [1:0] grant_store = 2'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [3:0] requests;
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$18 ) begin end
    grant = 2'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      2'h0:
        begin
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
        end
      2'h1:
        begin
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
        end
      2'h2:
        begin
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
        end
      2'h3:
        begin
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$18 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 2'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:454" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_north (clk, rst, inputs__0__valid, inputs__0__payload, inputs__1__valid, inputs__1__payload, inputs__2__valid, inputs__2__payload, inputs__3__valid, inputs__3__payload, input_ready, output__valid, output__payload, output__ready);
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  output [3:0] input_ready;
  wire [3:0] input_ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__0__payload;
  wire [79:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__1__payload;
  wire [79:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__2__payload;
  wire [79:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__3__payload;
  wire [79:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] output__payload;
  wire [75:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [77:0] \output__payload$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload$24.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$24.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload$24.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$26 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  assign \$1  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$2  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h9;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$2 , \$1  };
  assign input__0__valid = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$3 ;
  assign \$4  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$5  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h9;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$5 , \$4  };
  assign input__1__valid = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$6 ;
  assign \$7  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$8  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h9;
  assign \$9  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$8 , \$7  };
  assign input__2__valid = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$9 ;
  assign \$10  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$11  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'h9;
  assign \$12  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$11 , \$10  };
  assign input__3__valid = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:459" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_north.arbiter  arbiter (
    .clk(clk),
    .input__0__payload(input__0__payload),
    .input__0__ready(input__0__ready),
    .input__0__valid(input__0__valid),
    .input__1__payload(input__1__payload),
    .input__1__ready(input__1__ready),
    .input__1__valid(input__1__valid),
    .input__2__payload(input__2__payload),
    .input__2__ready(input__2__ready),
    .input__2__valid(input__2__valid),
    .input__3__payload(input__3__payload),
    .input__3__ready(input__3__ready),
    .input__3__valid(input__3__valid),
    .output__payload(\output__payload$24 ),
    .output__ready(output__ready),
    .output__valid(output__valid),
    .rst(rst)
  );
  assign \output__valid$22  = output__valid;
  assign \output__ready$26  = output__ready;
  assign output__payload = \output__payload$24 [75:0];
  assign \inputs__0__payload.last  = inputs__0__payload[75];
  assign \inputs__0__payload.target  = inputs__0__payload[79:76];
  assign \inputs__0__payload.target.port  = inputs__0__payload[78:76];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \inputs__1__payload.last  = inputs__1__payload[75];
  assign \inputs__1__payload.target  = inputs__1__payload[79:76];
  assign \inputs__1__payload.target.port  = inputs__1__payload[78:76];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \inputs__2__payload.last  = inputs__2__payload[75];
  assign \inputs__2__payload.target  = inputs__2__payload[79:76];
  assign \inputs__2__payload.target.port  = inputs__2__payload[78:76];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[79];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \inputs__3__payload.last  = inputs__3__payload[75];
  assign \inputs__3__payload.target  = inputs__3__payload[79:76];
  assign \inputs__3__payload.target.port  = inputs__3__payload[78:76];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[79];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign \output__payload.vc  = \output__payload$24 [75];
  assign \output__payload$24.p  = \output__payload$24 [75:0];
  assign \output__payload$24.p.vc  = \output__payload$24 [75];
  assign \output__payload$24.src  = \output__payload$24 [77:76];
  assign input__3__payload[75] = inputs__3__payload[79];
  assign input__3__payload[74:0] = inputs__3__payload[74:0];
  assign input__2__payload[75] = inputs__2__payload[79];
  assign input__2__payload[74:0] = inputs__2__payload[74:0];
  assign input__1__payload[75] = inputs__1__payload[79];
  assign input__1__payload[74:0] = inputs__1__payload[74:0];
  assign input_ready[3] = input__3__ready;
  assign input_ready[2] = input__2__ready;
  assign input_ready[1] = input__1__ready;
  assign input_ready[0] = input__0__ready;
  assign input__0__payload[75] = inputs__0__payload[79];
  assign input__0__payload[74:0] = inputs__0__payload[74:0];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_north.arbiter (clk, rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__0__payload, input__1__payload, input__2__payload, input__3__payload, output__valid, output__payload, input__0__ready, input__1__ready, input__2__ready, input__3__ready, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$19  = 0;
  reg \$1 ;
  reg [75:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [1:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg [1:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__0__payload;
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__1__payload;
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__2__payload;
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__3__payload;
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [77:0] output__payload;
  reg [77:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_north.arbiter.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$1  = input__0__valid;
      2'h1:
          \$1  = input__1__valid;
      2'h2:
          \$1  = input__2__valid;
      2'h3:
          \$1  = input__3__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$2  = input__0__payload;
      2'h1:
          \$2  = input__1__payload;
      2'h2:
          \$2  = input__2__payload;
      2'h3:
          \$2  = input__3__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    output__payload = 78'h00000000000000000000;
    if (transfer) begin
      output__payload[75:0] = \$2 ;
      output__payload[77:76] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            /* empty */;
        2'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    granted = 2'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$19 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[75:0];
  assign \output__payload.p.vc  = output__payload[75];
  assign \output__payload.src  = output__payload[77:76];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_north.arbiter.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$20  = 0;
  reg [1:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [1:0] grant;
  reg [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [1:0] grant_store;
  reg [1:0] grant_store = 2'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [3:0] requests;
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$20 ) begin end
    grant = 2'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      2'h0:
        begin
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
        end
      2'h1:
        begin
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
        end
      2'h2:
        begin
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
        end
      2'h3:
        begin
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$20 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 2'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:454" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_south (clk, rst, inputs__0__valid, inputs__0__payload, inputs__1__valid, inputs__1__payload, inputs__2__valid, inputs__2__payload, inputs__3__valid, inputs__3__payload, input_ready, output__valid, output__payload, output__ready);
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  output [3:0] input_ready;
  wire [3:0] input_ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__0__payload;
  wire [79:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__1__payload;
  wire [79:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__2__payload;
  wire [79:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__3__payload;
  wire [79:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] output__payload;
  wire [75:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [77:0] \output__payload$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload$24.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$24.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload$24.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$26 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  assign \$1  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h2;
  assign \$2  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'ha;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$2 , \$1  };
  assign input__0__valid = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$3 ;
  assign \$4  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h2;
  assign \$5  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'ha;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$5 , \$4  };
  assign input__1__valid = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$6 ;
  assign \$7  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h2;
  assign \$8  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'ha;
  assign \$9  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$8 , \$7  };
  assign input__2__valid = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$9 ;
  assign \$10  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h2;
  assign \$11  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'ha;
  assign \$12  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$11 , \$10  };
  assign input__3__valid = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:459" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_south.arbiter  arbiter (
    .clk(clk),
    .input__0__payload(input__0__payload),
    .input__0__ready(input__0__ready),
    .input__0__valid(input__0__valid),
    .input__1__payload(input__1__payload),
    .input__1__ready(input__1__ready),
    .input__1__valid(input__1__valid),
    .input__2__payload(input__2__payload),
    .input__2__ready(input__2__ready),
    .input__2__valid(input__2__valid),
    .input__3__payload(input__3__payload),
    .input__3__ready(input__3__ready),
    .input__3__valid(input__3__valid),
    .output__payload(\output__payload$24 ),
    .output__ready(output__ready),
    .output__valid(output__valid),
    .rst(rst)
  );
  assign \output__valid$22  = output__valid;
  assign \output__ready$26  = output__ready;
  assign output__payload = \output__payload$24 [75:0];
  assign \inputs__0__payload.last  = inputs__0__payload[75];
  assign \inputs__0__payload.target  = inputs__0__payload[79:76];
  assign \inputs__0__payload.target.port  = inputs__0__payload[78:76];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \inputs__1__payload.last  = inputs__1__payload[75];
  assign \inputs__1__payload.target  = inputs__1__payload[79:76];
  assign \inputs__1__payload.target.port  = inputs__1__payload[78:76];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \inputs__2__payload.last  = inputs__2__payload[75];
  assign \inputs__2__payload.target  = inputs__2__payload[79:76];
  assign \inputs__2__payload.target.port  = inputs__2__payload[78:76];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[79];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \inputs__3__payload.last  = inputs__3__payload[75];
  assign \inputs__3__payload.target  = inputs__3__payload[79:76];
  assign \inputs__3__payload.target.port  = inputs__3__payload[78:76];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[79];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign \output__payload.vc  = \output__payload$24 [75];
  assign \output__payload$24.p  = \output__payload$24 [75:0];
  assign \output__payload$24.p.vc  = \output__payload$24 [75];
  assign \output__payload$24.src  = \output__payload$24 [77:76];
  assign input__3__payload[75] = inputs__3__payload[79];
  assign input__3__payload[74:0] = inputs__3__payload[74:0];
  assign input__2__payload[75] = inputs__2__payload[79];
  assign input__2__payload[74:0] = inputs__2__payload[74:0];
  assign input__1__payload[75] = inputs__1__payload[79];
  assign input__1__payload[74:0] = inputs__1__payload[74:0];
  assign input_ready[3] = input__3__ready;
  assign input_ready[2] = input__2__ready;
  assign input_ready[1] = input__1__ready;
  assign input_ready[0] = input__0__ready;
  assign input__0__payload[75] = inputs__0__payload[79];
  assign input__0__payload[74:0] = inputs__0__payload[74:0];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_south.arbiter (clk, rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__0__payload, input__1__payload, input__2__payload, input__3__payload, output__valid, output__payload, input__0__ready, input__1__ready, input__2__ready, input__3__ready, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$21  = 0;
  reg \$1 ;
  reg [75:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [1:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg [1:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__0__payload;
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__1__payload;
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__2__payload;
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__3__payload;
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [77:0] output__payload;
  reg [77:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_south.arbiter.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$1  = input__0__valid;
      2'h1:
          \$1  = input__1__valid;
      2'h2:
          \$1  = input__2__valid;
      2'h3:
          \$1  = input__3__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$2  = input__0__payload;
      2'h1:
          \$2  = input__1__payload;
      2'h2:
          \$2  = input__2__payload;
      2'h3:
          \$2  = input__3__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    output__payload = 78'h00000000000000000000;
    if (transfer) begin
      output__payload[75:0] = \$2 ;
      output__payload[77:76] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            /* empty */;
        2'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    granted = 2'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$21 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[75:0];
  assign \output__payload.p.vc  = output__payload[75];
  assign \output__payload.src  = output__payload[77:76];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_south.arbiter.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$22  = 0;
  reg [1:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [1:0] grant;
  reg [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [1:0] grant_store;
  reg [1:0] grant_store = 2'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [3:0] requests;
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$22 ) begin end
    grant = 2'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      2'h0:
        begin
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
        end
      2'h1:
        begin
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
        end
      2'h2:
        begin
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
        end
      2'h3:
        begin
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$22 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 2'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:454" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_west (clk, rst, inputs__0__valid, inputs__0__payload, inputs__1__valid, inputs__1__payload, inputs__2__valid, inputs__2__payload, inputs__3__valid, inputs__3__payload, input_ready, output__valid, output__payload, output__ready);
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:447" *)
  output [3:0] input_ready;
  wire [3:0] input_ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__0__payload;
  wire [79:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__1__payload;
  wire [79:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__2__payload;
  wire [79:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] inputs__3__payload;
  wire [79:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  output [75:0] output__payload;
  wire [75:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [77:0] \output__payload$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload$24.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload$24.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload$24.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:444" *)
  wire \output__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$26 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  assign \$1  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 3'h4;
  assign \$2  = inputs__0__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hc;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$2 , \$1  };
  assign input__0__valid = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$3 ;
  assign \$4  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 3'h4;
  assign \$5  = inputs__1__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hc;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$5 , \$4  };
  assign input__1__valid = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$6 ;
  assign \$7  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 3'h4;
  assign \$8  = inputs__2__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hc;
  assign \$9  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$8 , \$7  };
  assign input__2__valid = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$9 ;
  assign \$10  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 3'h4;
  assign \$11  = inputs__3__payload[79:76] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 4'hc;
  assign \$12  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$11 , \$10  };
  assign input__3__valid = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:462" *) \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:459" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_west.arbiter  arbiter (
    .clk(clk),
    .input__0__payload(input__0__payload),
    .input__0__ready(input__0__ready),
    .input__0__valid(input__0__valid),
    .input__1__payload(input__1__payload),
    .input__1__ready(input__1__ready),
    .input__1__valid(input__1__valid),
    .input__2__payload(input__2__payload),
    .input__2__ready(input__2__ready),
    .input__2__valid(input__2__valid),
    .input__3__payload(input__3__payload),
    .input__3__ready(input__3__ready),
    .input__3__valid(input__3__valid),
    .output__payload(\output__payload$24 ),
    .output__ready(output__ready),
    .output__valid(output__valid),
    .rst(rst)
  );
  assign \output__valid$22  = output__valid;
  assign \output__ready$26  = output__ready;
  assign output__payload = \output__payload$24 [75:0];
  assign \inputs__0__payload.last  = inputs__0__payload[75];
  assign \inputs__0__payload.target  = inputs__0__payload[79:76];
  assign \inputs__0__payload.target.port  = inputs__0__payload[78:76];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[79];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \inputs__1__payload.last  = inputs__1__payload[75];
  assign \inputs__1__payload.target  = inputs__1__payload[79:76];
  assign \inputs__1__payload.target.port  = inputs__1__payload[78:76];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[79];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \inputs__2__payload.last  = inputs__2__payload[75];
  assign \inputs__2__payload.target  = inputs__2__payload[79:76];
  assign \inputs__2__payload.target.port  = inputs__2__payload[78:76];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[79];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \inputs__3__payload.last  = inputs__3__payload[75];
  assign \inputs__3__payload.target  = inputs__3__payload[79:76];
  assign \inputs__3__payload.target.port  = inputs__3__payload[78:76];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[79];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign \output__payload.vc  = \output__payload$24 [75];
  assign \output__payload$24.p  = \output__payload$24 [75:0];
  assign \output__payload$24.p.vc  = \output__payload$24 [75];
  assign \output__payload$24.src  = \output__payload$24 [77:76];
  assign input__3__payload[75] = inputs__3__payload[79];
  assign input__3__payload[74:0] = inputs__3__payload[74:0];
  assign input__2__payload[75] = inputs__2__payload[79];
  assign input__2__payload[74:0] = inputs__2__payload[74:0];
  assign input__1__payload[75] = inputs__1__payload[79];
  assign input__1__payload[74:0] = inputs__1__payload[74:0];
  assign input_ready[3] = input__3__ready;
  assign input_ready[2] = input__2__ready;
  assign input_ready[1] = input__1__ready;
  assign input_ready[0] = input__0__ready;
  assign input__0__payload[75] = inputs__0__payload[79];
  assign input__0__payload[74:0] = inputs__0__payload[74:0];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_west.arbiter (clk, rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__0__payload, input__1__payload, input__2__payload, input__3__payload, output__valid, output__payload, input__0__ready, input__1__ready, input__2__ready, input__3__ready, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$23  = 0;
  reg \$1 ;
  reg [75:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [1:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg [1:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__0__payload;
  wire [75:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__1__payload;
  wire [75:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__2__payload;
  wire [75:0] input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__2__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [75:0] input__3__payload;
  wire [75:0] input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__3__payload.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [77:0] output__payload;
  reg [77:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [75:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.vc ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [1:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_output_west.arbiter.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$1  = input__0__valid;
      2'h1:
          \$1  = input__1__valid;
      2'h2:
          \$1  = input__2__valid;
      2'h3:
          \$1  = input__3__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      2'h0:
          \$2  = input__0__payload;
      2'h1:
          \$2  = input__1__payload;
      2'h2:
          \$2  = input__2__payload;
      2'h3:
          \$2  = input__3__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    output__payload = 78'h00000000000000000000;
    if (transfer) begin
      output__payload[75:0] = \$2 ;
      output__payload[77:76] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        2'h0:
            /* empty */;
        2'h1:
            /* empty */;
        2'h2:
            /* empty */;
        2'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    granted = 2'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$23 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[75:0];
  assign \output__payload.p.vc  = output__payload[75];
  assign \output__payload.src  = output__payload[77:76];
  assign \input__0__payload.vc  = input__0__payload[75];
  assign \input__1__payload.vc  = input__1__payload[75];
  assign \input__2__payload.vc  = input__2__payload[75];
  assign \input__3__payload.vc  = input__3__payload[75];
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_output_west.arbiter.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$24  = 0;
  reg [1:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [1:0] grant;
  reg [1:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [1:0] grant_store;
  reg [1:0] grant_store = 2'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [3:0] requests;
  wire [3:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$24 ) begin end
    grant = 2'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      2'h0:
        begin
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
        end
      2'h1:
        begin
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
        end
      2'h2:
        begin
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
          if (requests[3]) begin
            grant = 2'h3;
          end
        end
      2'h3:
        begin
          if (requests[3]) begin
            grant = 2'h3;
          end
          if (requests[2]) begin
            grant = 2'h2;
          end
          if (requests[1]) begin
            grant = 2'h1;
          end
          if (requests[0]) begin
            grant = 2'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$24 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 2'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_south_arb (input__1__payload, clk, rst, input__0__valid, input__1__valid, output__ready, output__valid, output__payload, input__0__ready, input__1__ready, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$25  = 0;
  reg \$1 ;
  reg [79:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__0__payload;
  wire [79:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__1__payload;
  wire [79:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [80:0] output__payload;
  reg [80:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_south_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$1  = input__0__valid;
      1'h1:
          \$1  = input__1__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$2  = input__0__payload;
      1'h1:
          \$2  = input__1__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    output__payload = 81'h000000000000000000000;
    if (transfer) begin
      output__payload[79:0] = \$2 ;
      output__payload[80] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        1'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        1'h0:
            /* empty */;
        1'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    granted = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$25 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[79:0];
  assign \output__payload.p.last  = output__payload[75];
  assign \output__payload.p.target  = output__payload[79:76];
  assign \output__payload.p.target.port  = output__payload[78:76];
  assign \output__payload.p.target.vc_id  = output__payload[79];
  assign \output__payload.src  = output__payload[80];
  assign \input__0__payload.last  = input__0__payload[75];
  assign \input__0__payload.target  = input__0__payload[79:76];
  assign \input__0__payload.target.port  = input__0__payload[78:76];
  assign \input__0__payload.target.vc_id  = input__0__payload[79];
  assign \input__1__payload.last  = input__1__payload[75];
  assign \input__1__payload.target  = input__1__payload[79:76];
  assign \input__1__payload.target.port  = input__1__payload[78:76];
  assign \input__1__payload.target.vc_id  = input__1__payload[79];
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_south_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$26  = 0;
  reg \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output grant;
  reg grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output grant_store;
  reg grant_store = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [1:0] requests;
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$26 ) begin end
    grant = 1'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      1'h0:
        begin
          if (requests[0]) begin
            grant = 1'h0;
          end
          if (requests[1]) begin
            grant = 1'h1;
          end
        end
      1'h1:
        begin
          if (requests[1]) begin
            grant = 1'h1;
          end
          if (requests[0]) begin
            grant = 1'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$26 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 1'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_south_vc_0_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$27  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$27 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$27 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_south_vc_1_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$28  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$28 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$28 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_west_arb (input__1__payload, clk, rst, input__0__valid, input__1__valid, output__ready, output__valid, output__payload, input__0__ready, input__1__ready, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$29  = 0;
  reg \$1 ;
  reg [79:0] \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  reg \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:946" *)
  reg granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__0__payload;
  wire [79:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [79:0] input__1__payload;
  wire [79:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \input__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \input__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \input__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  output [80:0] output__payload;
  reg [80:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [79:0] \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [3:0] \output__payload.p.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire [2:0] \output__payload.p.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.p.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:929" *)
  wire \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:947" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:960" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:966" *) output__ready;
  assign \$8  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:975" *) output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:976" *)
  always @(posedge clk)
    fsm_state <= \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:941" *)
  \memory_mapped_router.RouterCrossbar.crossbar_west_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$1  = input__0__valid;
      1'h1:
          \$1  = input__1__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      1'h0:
          \$2  = input__0__payload;
      1'h1:
          \$2  = input__1__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    output__payload = 81'h000000000000000000000;
    if (transfer) begin
      output__payload[79:0] = \$2 ;
      output__payload[80] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        1'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        1'h0:
            /* empty */;
        1'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    granted = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$29 ) begin end
    \$9  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$7 ) begin
              \$9  = 1'h0;
            end else begin
              \$9  = 1'h1;
            end
          end
      1'h1:
          if (\$8 ) begin
            \$9  = 1'h0;
          end
    endcase
    if (rst) begin
      \$9  = 1'h0;
    end
  end
  assign \output__payload.p  = output__payload[79:0];
  assign \output__payload.p.last  = output__payload[75];
  assign \output__payload.p.target  = output__payload[79:76];
  assign \output__payload.p.target.port  = output__payload[78:76];
  assign \output__payload.p.target.vc_id  = output__payload[79];
  assign \output__payload.src  = output__payload[80];
  assign \input__0__payload.last  = input__0__payload[75];
  assign \input__0__payload.target  = input__0__payload[79:76];
  assign \input__0__payload.target.port  = input__0__payload[78:76];
  assign \input__0__payload.target.vc_id  = input__0__payload[79];
  assign \input__1__payload.last  = input__1__payload[75];
  assign \input__1__payload.target  = input__1__payload[79:76];
  assign \input__1__payload.target.port  = input__1__payload[78:76];
  assign \input__1__payload.target.vc_id  = input__1__payload[79];
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_west_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$30  = 0;
  reg \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output grant;
  reg grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output grant_store;
  reg grant_store = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [1:0] requests;
  wire [1:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$30 ) begin end
    grant = 1'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      1'h0:
        begin
          if (requests[0]) begin
            grant = 1'h0;
          end
          if (requests[1]) begin
            grant = 1'h1;
          end
        end
      1'h1:
        begin
          if (requests[1]) begin
            grant = 1'h1;
          end
          if (requests[0]) begin
            grant = 1'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$30 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 1'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_west_vc_0_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$31  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$31 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$31 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:484" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.crossbar_west_vc_1_tee (clk, rst, output__1__ready, output__0__ready, input__ready, output__0__valid, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$32  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  reg [1:0] \$12 ;
  reg \$13 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  reg in_stalled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:489" *)
  wire [1:0] next_stalled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [-1:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  reg [1:0] stalled = 2'h0;
  assign \$2  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:493" *) \$1 ;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) next_stalled;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:492" *) \$3 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__0__ready;
  assign \$5  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$4 ;
  assign \$6  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$6 ;
  assign output__0__valid = \$7  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[0];
  assign \$8  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) output__1__ready;
  assign \$9  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:496" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) in_stalled;
  assign \$11  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:487" *) \$10 ;
  assign output__1__valid = \$11  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:498" *) stalled[1];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:488" *)
  always @(posedge clk)
    stalled <= \$12 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:486" *)
  always @(posedge clk)
    in_stalled <= \$13 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$32 ) begin end
    \$12  = next_stalled;
    if (rst) begin
      \$12  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$32 ) begin end
    \$13  = \$2 ;
    if (rst) begin
      \$13  = 1'h0;
    end
  end
  assign next_stalled[1] = \$9 ;
  assign next_stalled[0] = \$5 ;
  assign \$1  = \$3 ;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:371" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator (credit_in__valid, \credit_in__payload$354 , \credit_in__valid$356 , \credit_in__payload$368 , \credit_in__valid$370 , \credit_in__payload$382 , \credit_in__valid$384 , clk, rst, outputs__0__ready, outputs__1__ready, outputs__2__ready, outputs__3__ready, outputs__4__ready, outputs__5__ready, outputs__6__ready, outputs__7__ready, outputs__8__ready, outputs__9__ready, inputs__0__ready, inputs__1__ready
, inputs__2__ready, inputs__3__ready, inputs__4__ready, inputs__5__ready, inputs__6__ready, inputs__7__ready, inputs__8__ready, inputs__9__ready, outputs__0__valid, outputs__1__valid, outputs__2__valid, outputs__3__valid, outputs__4__valid, outputs__5__valid, outputs__6__valid, outputs__7__valid, outputs__8__valid, outputs__9__valid, inputs__0__valid, inputs__1__valid, inputs__2__valid
, inputs__3__valid, inputs__4__valid, inputs__5__valid, inputs__6__valid, inputs__7__valid, inputs__8__valid, inputs__9__valid, inputs__0__payload, inputs__1__payload, inputs__2__payload, inputs__3__payload, inputs__4__payload, inputs__5__payload, inputs__6__payload, inputs__7__payload, inputs__8__payload, inputs__9__payload, credit_in__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$33  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$100 ;
  wire \$101 ;
  wire \$102 ;
  wire \$103 ;
  wire \$104 ;
  wire \$105 ;
  wire \$106 ;
  wire \$107 ;
  wire \$108 ;
  wire \$109 ;
  wire \$11 ;
  wire \$110 ;
  wire \$111 ;
  wire \$112 ;
  wire \$113 ;
  wire \$114 ;
  wire \$115 ;
  wire \$116 ;
  wire \$117 ;
  wire \$118 ;
  wire \$119 ;
  wire \$12 ;
  wire \$120 ;
  wire \$121 ;
  wire \$122 ;
  wire \$123 ;
  wire \$124 ;
  wire \$125 ;
  wire \$126 ;
  wire \$127 ;
  wire \$128 ;
  wire \$129 ;
  wire \$13 ;
  wire \$130 ;
  wire \$131 ;
  wire \$132 ;
  wire \$133 ;
  wire \$134 ;
  wire \$135 ;
  wire \$136 ;
  wire \$137 ;
  wire \$138 ;
  wire \$139 ;
  wire \$14 ;
  wire \$140 ;
  wire \$141 ;
  wire \$142 ;
  wire \$143 ;
  wire \$144 ;
  wire \$145 ;
  wire \$146 ;
  wire \$147 ;
  wire \$148 ;
  wire \$149 ;
  wire \$15 ;
  wire \$150 ;
  wire \$151 ;
  wire \$152 ;
  wire \$153 ;
  wire \$154 ;
  wire \$155 ;
  wire \$156 ;
  wire \$157 ;
  wire \$158 ;
  wire \$159 ;
  wire \$16 ;
  wire \$160 ;
  wire \$161 ;
  wire \$162 ;
  wire \$163 ;
  wire \$164 ;
  wire \$165 ;
  wire \$166 ;
  wire \$167 ;
  wire \$168 ;
  wire \$169 ;
  wire \$17 ;
  wire \$170 ;
  wire \$171 ;
  wire \$172 ;
  wire \$173 ;
  wire \$174 ;
  wire \$175 ;
  wire \$176 ;
  wire \$177 ;
  wire \$178 ;
  wire \$179 ;
  wire \$18 ;
  wire \$180 ;
  wire \$181 ;
  wire \$182 ;
  wire \$183 ;
  wire \$184 ;
  wire \$185 ;
  wire \$186 ;
  wire \$187 ;
  wire \$188 ;
  wire \$189 ;
  wire \$19 ;
  wire \$190 ;
  wire \$191 ;
  wire \$192 ;
  wire \$193 ;
  wire \$194 ;
  wire \$195 ;
  wire \$196 ;
  wire \$197 ;
  wire \$198 ;
  wire \$199 ;
  wire \$2 ;
  wire \$20 ;
  wire \$200 ;
  wire \$201 ;
  wire \$202 ;
  wire \$203 ;
  wire \$204 ;
  wire \$205 ;
  wire \$206 ;
  wire \$207 ;
  wire \$208 ;
  wire \$209 ;
  wire \$21 ;
  wire \$210 ;
  wire \$211 ;
  wire \$212 ;
  wire \$213 ;
  wire \$214 ;
  wire \$215 ;
  wire \$216 ;
  wire \$217 ;
  wire \$218 ;
  wire \$219 ;
  wire \$22 ;
  wire \$220 ;
  wire \$221 ;
  wire \$222 ;
  wire \$223 ;
  wire \$224 ;
  wire \$225 ;
  wire \$226 ;
  wire \$227 ;
  wire \$228 ;
  wire \$229 ;
  wire \$23 ;
  wire \$230 ;
  wire \$231 ;
  wire \$232 ;
  wire \$233 ;
  wire \$234 ;
  wire \$235 ;
  wire \$236 ;
  wire \$237 ;
  wire \$238 ;
  wire \$239 ;
  wire \$24 ;
  wire \$240 ;
  wire \$241 ;
  wire \$242 ;
  wire \$243 ;
  wire \$244 ;
  wire \$245 ;
  wire \$246 ;
  wire \$247 ;
  wire \$248 ;
  wire \$249 ;
  wire \$25 ;
  wire \$250 ;
  wire \$251 ;
  wire \$252 ;
  wire \$253 ;
  wire \$254 ;
  wire \$255 ;
  wire \$256 ;
  wire \$257 ;
  wire \$258 ;
  wire \$259 ;
  wire \$26 ;
  wire \$260 ;
  wire \$261 ;
  wire \$262 ;
  wire \$263 ;
  wire \$264 ;
  wire \$265 ;
  wire \$266 ;
  wire \$267 ;
  wire \$268 ;
  wire \$269 ;
  wire \$27 ;
  wire \$270 ;
  wire \$271 ;
  wire \$272 ;
  wire \$273 ;
  wire \$274 ;
  wire \$275 ;
  wire \$276 ;
  wire \$277 ;
  wire \$278 ;
  wire \$279 ;
  wire \$28 ;
  wire \$280 ;
  wire \$281 ;
  wire \$282 ;
  wire \$283 ;
  wire \$284 ;
  wire \$285 ;
  wire \$286 ;
  wire \$287 ;
  wire \$288 ;
  wire \$289 ;
  wire \$29 ;
  wire \$290 ;
  wire \$291 ;
  wire \$292 ;
  wire \$293 ;
  wire \$294 ;
  wire \$295 ;
  wire \$296 ;
  wire \$297 ;
  wire \$298 ;
  wire \$299 ;
  wire \$3 ;
  wire \$30 ;
  wire \$300 ;
  wire \$301 ;
  wire \$302 ;
  wire \$303 ;
  wire \$304 ;
  wire \$305 ;
  wire \$306 ;
  wire \$307 ;
  wire \$308 ;
  wire \$309 ;
  wire \$31 ;
  wire \$310 ;
  wire \$311 ;
  wire \$312 ;
  wire \$313 ;
  wire \$314 ;
  wire \$315 ;
  wire \$316 ;
  wire \$317 ;
  wire \$318 ;
  wire \$319 ;
  wire \$32 ;
  wire \$320 ;
  wire \$321 ;
  wire \$322 ;
  wire \$33 ;
  wire \$34 ;
  wire \$35 ;
  wire \$36 ;
  wire \$37 ;
  wire \$38 ;
  wire \$39 ;
  wire \$4 ;
  wire \$40 ;
  wire \$41 ;
  wire \$42 ;
  wire \$43 ;
  wire \$44 ;
  wire \$45 ;
  wire \$46 ;
  wire \$47 ;
  wire \$48 ;
  wire \$49 ;
  wire \$5 ;
  wire \$50 ;
  wire \$51 ;
  wire \$52 ;
  wire \$53 ;
  wire \$54 ;
  wire \$55 ;
  wire \$56 ;
  wire \$57 ;
  wire \$58 ;
  wire \$59 ;
  wire \$6 ;
  wire \$60 ;
  wire \$61 ;
  wire \$62 ;
  wire \$63 ;
  wire \$64 ;
  wire \$65 ;
  wire \$66 ;
  wire \$67 ;
  wire \$68 ;
  wire \$69 ;
  wire \$7 ;
  wire \$70 ;
  wire \$71 ;
  wire \$72 ;
  reg [2:0] \$73 ;
  wire \$74 ;
  wire \$75 ;
  wire \$76 ;
  wire \$77 ;
  wire \$78 ;
  wire \$79 ;
  wire \$8 ;
  wire \$80 ;
  wire \$81 ;
  reg [2:0] \$82 ;
  wire \$83 ;
  wire \$84 ;
  wire \$85 ;
  wire \$86 ;
  wire \$87 ;
  wire \$88 ;
  wire \$89 ;
  wire \$9 ;
  wire \$90 ;
  wire \$91 ;
  wire \$92 ;
  wire \$93 ;
  wire \$94 ;
  wire \$95 ;
  wire \$96 ;
  wire \$97 ;
  wire \$98 ;
  wire \$99 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload$104 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload$126 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload$148 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload$170 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload$192 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \$signature__payload$214 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \$signature__payload$236 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload$56 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  reg [3:0] \$signature__payload$82 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$107 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$129 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$151 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$173 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$195 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$217 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$239 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$59 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \$signature__ready$85 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$102 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$124 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$146 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$168 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$190 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$212 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$234 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$54 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \$signature__valid$80 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] credit__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__0__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__0__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire credit__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] credit__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__1__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__1__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire credit__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] credit__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__2__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__2__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire credit__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [11:0] credit__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__3__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [5:0] \credit__3__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire credit__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] credit_in__payload;
  wire [11:0] credit_in__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] \credit_in__payload$354 ;
  wire [11:0] \credit_in__payload$354 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload$354[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload$354[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] \credit_in__payload$368 ;
  wire [11:0] \credit_in__payload$368 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload$368[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload$368[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [11:0] \credit_in__payload$382 ;
  wire [11:0] \credit_in__payload$382 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload$382[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload$382[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit_in__valid;
  wire credit_in__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input \credit_in__valid$356 ;
  wire \credit_in__valid$356 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input \credit_in__valid$370 ;
  wire \credit_in__valid$370 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input \credit_in__valid$384 ;
  wire \credit_in__valid$384 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$109 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$131 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$153 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$175 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$197 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$219 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__0__payload$344 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__0__payload$358 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__0__payload$372 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__0__payload$386 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$39 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$63 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__0__payload$87 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$242 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$243 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$244 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$245 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$246 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$247 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$248 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$259 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$260 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$345 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$359 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$373 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__0__ready$387 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$108 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$130 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$152 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$174 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$196 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$218 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$346 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$360 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$374 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$38 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$388 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$60 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__0__valid$86 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$111 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$133 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$155 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$177 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$199 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$221 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__1__payload$349 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__1__payload$363 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__1__payload$377 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \input__1__payload$391 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$41 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$67 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__1__payload$89 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$251 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$252 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$253 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$254 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$255 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$256 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$257 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$268 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$269 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$350 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$364 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$378 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__1__ready$392 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$110 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$132 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$154 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$176 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$198 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$220 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$351 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$365 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$379 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$393 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$40 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$64 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__1__valid$88 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$113 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$135 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$157 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$179 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$201 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$223 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$43 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$69 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__2__payload$91 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$262 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$263 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$264 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$265 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$266 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$277 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$278 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$279 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__2__ready$280 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$112 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$134 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$156 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$178 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$200 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$222 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$42 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$68 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__2__valid$90 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$115 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$137 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$159 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$181 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$203 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$225 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$45 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$71 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__3__payload$93 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$271 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$272 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$273 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$274 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$275 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$286 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$287 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$288 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__3__ready$289 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$114 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$136 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$158 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$180 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$202 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$224 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$44 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$70 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__3__valid$92 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$117 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$139 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$161 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$183 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$205 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$227 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$47 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$73 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__4__payload$95 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$282 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$283 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$284 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$295 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$296 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$297 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$298 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$299 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__4__ready$300 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$116 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$138 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$160 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$182 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$204 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$226 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$46 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$72 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__4__valid$94 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$119 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$141 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$163 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$185 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$207 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$229 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$49 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$75 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__5__payload$97 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$291 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$292 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$293 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$304 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$305 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$306 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$307 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$308 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__5__ready$309 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$118 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$140 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$162 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$184 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$206 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$228 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$48 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$74 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__5__valid$96 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$121 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$143 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$165 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$187 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$209 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$231 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$51 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$77 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__6__payload$99 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$302 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$313 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$314 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$315 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$316 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$317 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$318 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$319 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__6__ready$320 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$120 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$142 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$164 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$186 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$208 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$230 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$50 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$76 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__6__valid$98 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$101 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$123 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$145 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$167 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$189 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$211 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$233 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$53 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire \input__7__payload$79 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$311 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$322 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$323 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$324 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$325 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$326 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$327 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$328 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \input__7__ready$329 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$100 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$122 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$144 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$166 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$188 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$210 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$232 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$52 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \input__7__valid$78 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__0__payload;
  wire [4:0] inputs__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__0__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__0__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__0__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__0__ready;
  wire inputs__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__0__valid;
  wire inputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__1__payload;
  wire [4:0] inputs__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__1__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__1__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__1__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__1__ready;
  wire inputs__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__1__valid;
  wire inputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__2__payload;
  wire [4:0] inputs__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__2__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__2__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__2__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__2__ready;
  wire inputs__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__2__valid;
  wire inputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__3__payload;
  wire [4:0] inputs__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__3__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__3__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__3__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__3__ready;
  wire inputs__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__3__valid;
  wire inputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__4__payload;
  wire [4:0] inputs__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__4__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__4__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__4__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__4__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__4__ready;
  wire inputs__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__4__valid;
  wire inputs__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__5__payload;
  wire [4:0] inputs__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__5__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__5__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__5__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__5__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__5__ready;
  wire inputs__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__5__valid;
  wire inputs__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__6__payload;
  wire [4:0] inputs__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__6__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__6__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__6__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__6__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__6__ready;
  wire inputs__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__6__valid;
  wire inputs__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__7__payload;
  wire [4:0] inputs__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__7__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__7__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__7__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__7__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__7__ready;
  wire inputs__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__7__valid;
  wire inputs__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__8__payload;
  wire [4:0] inputs__8__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__8__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__8__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__8__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__8__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__8__ready;
  wire inputs__8__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__8__valid;
  wire inputs__8__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  input [4:0] inputs__9__payload;
  wire [4:0] inputs__9__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__9__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [3:0] \inputs__9__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire [2:0] \inputs__9__payload.target.port ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1702" *)
  wire \inputs__9__payload.target.vc_id ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output inputs__9__ready;
  wire inputs__9__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input inputs__9__valid;
  wire inputs__9__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \output__0__payload$362 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \output__0__payload$376 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \output__0__payload$390 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg \output__0__ready$361 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg \output__0__ready$375 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg \output__0__ready$389 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$399 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$401 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__0__valid$403 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \output__1__payload$367 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \output__1__payload$381 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] \output__1__payload$395 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg \output__1__ready$366 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg \output__1__ready$380 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg \output__1__ready$394 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$400 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$402 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__1__valid$404 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$105 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$105.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$105.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$127 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$127.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$127.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$149 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$149.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$149.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$171 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$171.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$171.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$193 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$193.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$193.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$215 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$215.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$215.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$237 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$237.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$237.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$57 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$57.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$57.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [3:0] \output__payload$83 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload$83.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload$83.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$106 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$128 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$150 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$172 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$194 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$216 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$238 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  reg \output__ready$58 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \output__ready$84 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$103 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$125 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$147 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$169 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$191 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$213 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$235 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$55 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \output__valid$81 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__0__ready;
  wire outputs__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__0__valid;
  wire outputs__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__1__ready;
  wire outputs__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__1__valid;
  wire outputs__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__2__ready;
  wire outputs__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__2__valid;
  wire outputs__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__3__ready;
  wire outputs__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__3__valid;
  wire outputs__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__4__ready;
  wire outputs__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__4__valid;
  wire outputs__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__5__ready;
  wire outputs__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__5__valid;
  wire outputs__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__6__ready;
  wire outputs__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__6__valid;
  wire outputs__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__7__ready;
  wire outputs__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__7__valid;
  wire outputs__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__8__ready;
  wire outputs__8__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__8__valid;
  wire outputs__8__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input outputs__9__ready;
  wire outputs__9__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output outputs__9__valid;
  wire outputs__9__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  assign \$1  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__2__payload[3:0];
  assign input__0__valid = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$1 ;
  assign \$2  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__3__payload[3:0];
  assign input__1__valid = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$2 ;
  assign \$3  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__4__payload[3:0];
  assign input__2__valid = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$3 ;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__5__payload[3:0];
  assign input__3__valid = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$4 ;
  assign \$5  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__6__payload[3:0];
  assign input__4__valid = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$5 ;
  assign \$6  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__7__payload[3:0];
  assign input__5__valid = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$6 ;
  assign \$7  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__8__payload[3:0];
  assign input__6__valid = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$7 ;
  assign \$8  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) inputs__9__payload[3:0];
  assign input__7__valid = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$8 ;
  assign \$9  = inputs__2__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__0__valid$38  = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$9 ;
  assign \$10  = inputs__3__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__1__valid$40  = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$10 ;
  assign \$11  = inputs__4__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__2__valid$42  = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$11 ;
  assign \$12  = inputs__5__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__3__valid$44  = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$12 ;
  assign \$13  = inputs__6__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__4__valid$46  = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$13 ;
  assign \$14  = inputs__7__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__5__valid$48  = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$14 ;
  assign \$15  = inputs__8__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__6__valid$50  = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$15 ;
  assign \$16  = inputs__9__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h8;
  assign \input__7__valid$52  = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$16 ;
  assign \$17  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__0__valid$60  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$17 ;
  assign \$18  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__1__valid$64  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$18 ;
  assign \$19  = inputs__4__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__2__valid$68  = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$19 ;
  assign \$20  = inputs__5__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__3__valid$70  = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$20 ;
  assign \$21  = inputs__6__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__4__valid$72  = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$21 ;
  assign \$22  = inputs__7__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__5__valid$74  = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$22 ;
  assign \$23  = inputs__8__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__6__valid$76  = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$23 ;
  assign \$24  = inputs__9__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 1'h1;
  assign \input__7__valid$78  = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$24 ;
  assign \$25  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__0__valid$86  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$25 ;
  assign \$26  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__1__valid$88  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$26 ;
  assign \$27  = inputs__4__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__2__valid$90  = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$27 ;
  assign \$28  = inputs__5__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__3__valid$92  = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$28 ;
  assign \$29  = inputs__6__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__4__valid$94  = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$29 ;
  assign \$30  = inputs__7__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__5__valid$96  = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$30 ;
  assign \$31  = inputs__8__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__6__valid$98  = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$31 ;
  assign \$32  = inputs__9__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'h9;
  assign \input__7__valid$100  = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$32 ;
  assign \$33  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__0__valid$108  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$33 ;
  assign \$34  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__1__valid$110  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$34 ;
  assign \$35  = inputs__2__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__2__valid$112  = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$35 ;
  assign \$36  = inputs__3__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__3__valid$114  = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$36 ;
  assign \$37  = inputs__6__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__4__valid$116  = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$37 ;
  assign \$38  = inputs__7__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__5__valid$118  = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$38 ;
  assign \$39  = inputs__8__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__6__valid$120  = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$39 ;
  assign \$40  = inputs__9__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h2;
  assign \input__7__valid$122  = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$40 ;
  assign \$41  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__0__valid$130  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$41 ;
  assign \$42  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__1__valid$132  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$42 ;
  assign \$43  = inputs__2__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__2__valid$134  = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$43 ;
  assign \$44  = inputs__3__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__3__valid$136  = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$44 ;
  assign \$45  = inputs__6__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__4__valid$138  = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$45 ;
  assign \$46  = inputs__7__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__5__valid$140  = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$46 ;
  assign \$47  = inputs__8__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__6__valid$142  = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$47 ;
  assign \$48  = inputs__9__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'ha;
  assign \input__7__valid$144  = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$48 ;
  assign \$49  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__0__valid$152  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$49 ;
  assign \$50  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__1__valid$154  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$50 ;
  assign \$51  = inputs__2__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__2__valid$156  = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$51 ;
  assign \$52  = inputs__3__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__3__valid$158  = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$52 ;
  assign \$53  = inputs__4__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__4__valid$160  = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$53 ;
  assign \$54  = inputs__5__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__5__valid$162  = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$54 ;
  assign \$55  = inputs__8__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__6__valid$164  = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$55 ;
  assign \$56  = inputs__9__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 2'h3;
  assign \input__7__valid$166  = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$56 ;
  assign \$57  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__0__valid$174  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$57 ;
  assign \$58  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__1__valid$176  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$58 ;
  assign \$59  = inputs__2__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__2__valid$178  = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$59 ;
  assign \$60  = inputs__3__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__3__valid$180  = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$60 ;
  assign \$61  = inputs__4__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__4__valid$182  = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$61 ;
  assign \$62  = inputs__5__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__5__valid$184  = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$62 ;
  assign \$63  = inputs__8__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__6__valid$186  = inputs__8__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$63 ;
  assign \$64  = inputs__9__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hb;
  assign \input__7__valid$188  = inputs__9__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$64 ;
  assign \$65  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__0__valid$196  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$65 ;
  assign \$66  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__1__valid$198  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$66 ;
  assign \$67  = inputs__2__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__2__valid$200  = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$67 ;
  assign \$68  = inputs__3__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__3__valid$202  = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$68 ;
  assign \$69  = inputs__4__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__4__valid$204  = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$69 ;
  assign \$70  = inputs__5__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__5__valid$206  = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$70 ;
  assign \$71  = inputs__6__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__6__valid$208  = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$71 ;
  assign \$72  = inputs__7__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 3'h4;
  assign \input__7__valid$210  = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$72 ;
  assign \$74  = inputs__0__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__0__valid$218  = inputs__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$74 ;
  assign \$75  = inputs__1__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__1__valid$220  = inputs__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$75 ;
  assign \$76  = inputs__2__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__2__valid$222  = inputs__2__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$76 ;
  assign \$77  = inputs__3__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__3__valid$224  = inputs__3__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$77 ;
  assign \$78  = inputs__4__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__4__valid$226  = inputs__4__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$78 ;
  assign \$79  = inputs__5__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__5__valid$228  = inputs__5__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$79 ;
  assign \$80  = inputs__6__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__6__valid$230  = inputs__6__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$80 ;
  assign \$81  = inputs__7__payload[3:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/data.py:885" *) 4'hc;
  assign \input__7__valid$232  = inputs__7__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:391" *) \$81 ;
  assign \$83  = input__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$60 ;
  assign \$84  = \input__0__ready$242  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$86 ;
  assign \$85  = \input__0__ready$243  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$108 ;
  assign \$86  = \input__0__ready$244  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$130 ;
  assign \$87  = \input__0__ready$245  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$152 ;
  assign \$88  = \input__0__ready$246  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$174 ;
  assign \$89  = \input__0__ready$247  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$196 ;
  assign \$90  = \input__0__ready$248  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$218 ;
  assign inputs__0__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$90 , \$89 , \$88 , \$87 , \$86 , \$85 , \$84 , \$83  };
  assign \$91  = input__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$64 ;
  assign \$92  = \input__1__ready$251  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$88 ;
  assign \$93  = \input__1__ready$252  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$110 ;
  assign \$94  = \input__1__ready$253  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$132 ;
  assign \$95  = \input__1__ready$254  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$154 ;
  assign \$96  = \input__1__ready$255  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$176 ;
  assign \$97  = \input__1__ready$256  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$198 ;
  assign \$98  = \input__1__ready$257  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$220 ;
  assign inputs__1__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$98 , \$97 , \$96 , \$95 , \$94 , \$93 , \$92 , \$91  };
  assign \$99  = \input__0__ready$259  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__0__valid;
  assign \$100  = \input__0__ready$260  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__0__valid$38 ;
  assign \$101  = input__2__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$112 ;
  assign \$102  = \input__2__ready$262  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$134 ;
  assign \$103  = \input__2__ready$263  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$156 ;
  assign \$104  = \input__2__ready$264  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$178 ;
  assign \$105  = \input__2__ready$265  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$200 ;
  assign \$106  = \input__2__ready$266  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$222 ;
  assign inputs__2__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$106 , \$105 , \$104 , \$103 , \$102 , \$101 , \$100 , \$99  };
  assign \$107  = \input__1__ready$268  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__1__valid;
  assign \$108  = \input__1__ready$269  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__1__valid$40 ;
  assign \$109  = input__3__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$114 ;
  assign \$110  = \input__3__ready$271  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$136 ;
  assign \$111  = \input__3__ready$272  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$158 ;
  assign \$112  = \input__3__ready$273  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$180 ;
  assign \$113  = \input__3__ready$274  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$202 ;
  assign \$114  = \input__3__ready$275  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$224 ;
  assign inputs__3__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$114 , \$113 , \$112 , \$111 , \$110 , \$109 , \$108 , \$107  };
  assign \$115  = \input__2__ready$277  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__2__valid;
  assign \$116  = \input__2__ready$278  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$42 ;
  assign \$117  = \input__2__ready$279  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$68 ;
  assign \$118  = \input__2__ready$280  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__2__valid$90 ;
  assign \$119  = input__4__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$160 ;
  assign \$120  = \input__4__ready$282  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$182 ;
  assign \$121  = \input__4__ready$283  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$204 ;
  assign \$122  = \input__4__ready$284  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$226 ;
  assign inputs__4__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$122 , \$121 , \$120 , \$119 , \$118 , \$117 , \$116 , \$115  };
  assign \$123  = \input__3__ready$286  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__3__valid;
  assign \$124  = \input__3__ready$287  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$44 ;
  assign \$125  = \input__3__ready$288  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$70 ;
  assign \$126  = \input__3__ready$289  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__3__valid$92 ;
  assign \$127  = input__5__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$162 ;
  assign \$128  = \input__5__ready$291  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$184 ;
  assign \$129  = \input__5__ready$292  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$206 ;
  assign \$130  = \input__5__ready$293  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$228 ;
  assign inputs__5__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$130 , \$129 , \$128 , \$127 , \$126 , \$125 , \$124 , \$123  };
  assign \$131  = \input__4__ready$295  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__4__valid;
  assign \$132  = \input__4__ready$296  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$46 ;
  assign \$133  = \input__4__ready$297  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$72 ;
  assign \$134  = \input__4__ready$298  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$94 ;
  assign \$135  = \input__4__ready$299  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$116 ;
  assign \$136  = \input__4__ready$300  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__4__valid$138 ;
  assign \$137  = input__6__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$208 ;
  assign \$138  = \input__6__ready$302  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$230 ;
  assign inputs__6__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$138 , \$137 , \$136 , \$135 , \$134 , \$133 , \$132 , \$131  };
  assign \$139  = \input__5__ready$304  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__5__valid;
  assign \$140  = \input__5__ready$305  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$48 ;
  assign \$141  = \input__5__ready$306  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$74 ;
  assign \$142  = \input__5__ready$307  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$96 ;
  assign \$143  = \input__5__ready$308  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$118 ;
  assign \$144  = \input__5__ready$309  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__5__valid$140 ;
  assign \$145  = input__7__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$210 ;
  assign \$146  = \input__7__ready$311  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$232 ;
  assign inputs__7__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$146 , \$145 , \$144 , \$143 , \$142 , \$141 , \$140 , \$139  };
  assign \$147  = \input__6__ready$313  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__6__valid;
  assign \$148  = \input__6__ready$314  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$50 ;
  assign \$149  = \input__6__ready$315  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$76 ;
  assign \$150  = \input__6__ready$316  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$98 ;
  assign \$151  = \input__6__ready$317  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$120 ;
  assign \$152  = \input__6__ready$318  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$142 ;
  assign \$153  = \input__6__ready$319  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$164 ;
  assign \$154  = \input__6__ready$320  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__6__valid$186 ;
  assign inputs__8__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$154 , \$153 , \$152 , \$151 , \$150 , \$149 , \$148 , \$147  };
  assign \$155  = \input__7__ready$322  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) input__7__valid;
  assign \$156  = \input__7__ready$323  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$52 ;
  assign \$157  = \input__7__ready$324  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$78 ;
  assign \$158  = \input__7__ready$325  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$100 ;
  assign \$159  = \input__7__ready$326  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$122 ;
  assign \$160  = \input__7__ready$327  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$144 ;
  assign \$161  = \input__7__ready$328  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$166 ;
  assign \$162  = \input__7__ready$329  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:394" *) \input__7__valid$188 ;
  assign inputs__9__ready = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:403" *) { \$162 , \$161 , \$160 , \$159 , \$158 , \$157 , \$156 , \$155  };
  assign \$163  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$signature__payload$82 ;
  assign \$164  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$163 ;
  assign \$165  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$signature__payload$104 ;
  assign \$166  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$165 ;
  assign \$167  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$signature__payload$126 ;
  assign \$168  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$167 ;
  assign \$169  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$signature__payload$148 ;
  assign \$170  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$169 ;
  assign \$171  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$signature__payload$170 ;
  assign \$172  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$171 ;
  assign \$173  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$signature__payload$192 ;
  assign \$174  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$173 ;
  assign \$175  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$73 ;
  assign \$176  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$175 ;
  assign \$177  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$82 ;
  assign \$178  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$177 ;
  assign outputs__0__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$178 , \$176 , \$174 , \$172 , \$170 , \$168 , \$166 , \$164  };
  assign \$179  = \$signature__payload$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$180  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$179 ;
  assign \$181  = \$signature__payload$104  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$182  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$181 ;
  assign \$183  = \$signature__payload$126  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$184  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$183 ;
  assign \$185  = \$signature__payload$148  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$186  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$185 ;
  assign \$187  = \$signature__payload$170  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$188  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$187 ;
  assign \$189  = \$signature__payload$192  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$190  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$189 ;
  assign \$191  = \$73  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$192  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$191 ;
  assign \$193  = \$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 1'h1;
  assign \$194  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$193 ;
  assign outputs__1__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$194 , \$192 , \$190 , \$188 , \$186 , \$184 , \$182 , \$180  };
  assign \$195  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$196  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$195 ;
  assign \$197  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$198  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$197 ;
  assign \$199  = \$signature__payload$126  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$200  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$199 ;
  assign \$201  = \$signature__payload$148  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$202  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$201 ;
  assign \$203  = \$signature__payload$170  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$204  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$203 ;
  assign \$205  = \$signature__payload$192  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$206  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$205 ;
  assign \$207  = \$73  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$208  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$207 ;
  assign \$209  = \$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h2;
  assign \$210  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$209 ;
  assign outputs__2__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$210 , \$208 , \$206 , \$204 , \$202 , \$200 , \$198 , \$196  };
  assign \$211  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$212  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$211 ;
  assign \$213  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$214  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$213 ;
  assign \$215  = \$signature__payload$126  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$216  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$215 ;
  assign \$217  = \$signature__payload$148  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$218  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$217 ;
  assign \$219  = \$signature__payload$170  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$220  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$219 ;
  assign \$221  = \$signature__payload$192  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$222  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$221 ;
  assign \$223  = \$73  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$224  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$223 ;
  assign \$225  = \$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 2'h3;
  assign \$226  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$225 ;
  assign outputs__3__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$226 , \$224 , \$222 , \$220 , \$218 , \$216 , \$214 , \$212  };
  assign \$227  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$228  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$227 ;
  assign \$229  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$230  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$229 ;
  assign \$231  = \$signature__payload$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$232  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$231 ;
  assign \$233  = \$signature__payload$104  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$234  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$233 ;
  assign \$235  = \$signature__payload$170  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$236  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$235 ;
  assign \$237  = \$signature__payload$192  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$238  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$237 ;
  assign \$239  = \$73  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$240  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$239 ;
  assign \$241  = \$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h4;
  assign \$242  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$241 ;
  assign outputs__4__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$242 , \$240 , \$238 , \$236 , \$234 , \$232 , \$230 , \$228  };
  assign \$243  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$244  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$243 ;
  assign \$245  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$246  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$245 ;
  assign \$247  = \$signature__payload$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$248  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$247 ;
  assign \$249  = \$signature__payload$104  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$250  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$249 ;
  assign \$251  = \$signature__payload$170  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$252  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$251 ;
  assign \$253  = \$signature__payload$192  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$254  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$253 ;
  assign \$255  = \$73  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$256  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$255 ;
  assign \$257  = \$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h5;
  assign \$258  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$257 ;
  assign outputs__5__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$258 , \$256 , \$254 , \$252 , \$250 , \$248 , \$246 , \$244  };
  assign \$259  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$260  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$259 ;
  assign \$261  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$262  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$261 ;
  assign \$263  = \$signature__payload$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$264  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$263 ;
  assign \$265  = \$signature__payload$104  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$266  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$265 ;
  assign \$267  = \$signature__payload$126  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$268  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$267 ;
  assign \$269  = \$signature__payload$148  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$270  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$269 ;
  assign \$271  = \$73  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$272  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$271 ;
  assign \$273  = \$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h6;
  assign \$274  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$273 ;
  assign outputs__6__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$274 , \$272 , \$270 , \$268 , \$266 , \$264 , \$262 , \$260  };
  assign \$275  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$276  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$275 ;
  assign \$277  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$278  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$277 ;
  assign \$279  = \$signature__payload$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$280  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$279 ;
  assign \$281  = \$signature__payload$104  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$282  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$281 ;
  assign \$283  = \$signature__payload$126  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$284  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$283 ;
  assign \$285  = \$signature__payload$148  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$286  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$285 ;
  assign \$287  = \$73  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$288  = \output__0__valid$403  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$287 ;
  assign \$289  = \$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 3'h7;
  assign \$290  = \output__1__valid$404  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$289 ;
  assign outputs__7__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$290 , \$288 , \$286 , \$284 , \$282 , \$280 , \$278 , \$276  };
  assign \$291  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$292  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$291 ;
  assign \$293  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$294  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$293 ;
  assign \$295  = \$signature__payload$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$296  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$295 ;
  assign \$297  = \$signature__payload$104  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$298  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$297 ;
  assign \$299  = \$signature__payload$126  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$300  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$299 ;
  assign \$301  = \$signature__payload$148  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$302  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$301 ;
  assign \$303  = \$signature__payload$170  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$304  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$303 ;
  assign \$305  = \$signature__payload$192  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h8;
  assign \$306  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$305 ;
  assign outputs__8__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$306 , \$304 , \$302 , \$300 , \$298 , \$296 , \$294 , \$292  };
  assign \$307  = \$signature__payload  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$308  = \$signature__valid  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$307 ;
  assign \$309  = \$signature__payload$56  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$310  = \$signature__valid$54  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$309 ;
  assign \$311  = \$signature__payload$82  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$312  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$311 ;
  assign \$313  = \$signature__payload$104  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$314  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$313 ;
  assign \$315  = \$signature__payload$126  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$316  = \output__0__valid$399  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$315 ;
  assign \$317  = \$signature__payload$148  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$318  = \output__1__valid$400  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$317 ;
  assign \$319  = \$signature__payload$170  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$320  = \output__0__valid$401  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$319 ;
  assign \$321  = \$signature__payload$192  == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) 4'h9;
  assign \$322  = \output__1__valid$402  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:435" *) \$321 ;
  assign outputs__9__valid = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:438" *) { \$322 , \$320 , \$318 , \$316 , \$314 , \$312 , \$310 , \$308  };
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:409" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east  credit_counter_tx_east (
    .clk(clk),
    .credit_in__payload(\credit_in__payload$368 ),
    .credit_in__valid(\credit_in__valid$370 ),
    .input__0__ready(\output__ready$172 ),
    .input__0__valid(\$signature__valid$168 ),
    .input__1__ready(\output__ready$194 ),
    .input__1__valid(\$signature__valid$190 ),
    .output__0__payload(\$signature__payload$170 ),
    .output__0__ready(\output__0__ready$375 ),
    .output__0__valid(\output__0__valid$401 ),
    .output__1__payload(\$signature__payload$192 ),
    .output__1__ready(\output__1__ready$380 ),
    .output__1__valid(\output__1__valid$402 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_0_arb  credit_counter_tx_east_vc_0_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(\input__0__ready$245 ),
    .input__0__valid(\input__0__valid$152 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(\input__1__ready$254 ),
    .input__1__valid(\input__1__valid$154 ),
    .input__2__payload(inputs__2__payload[4]),
    .input__2__ready(\input__2__ready$263 ),
    .input__2__valid(\input__2__valid$156 ),
    .input__3__payload(inputs__3__payload[4]),
    .input__3__ready(\input__3__ready$272 ),
    .input__3__valid(\input__3__valid$158 ),
    .input__4__payload(inputs__4__payload[4]),
    .input__4__ready(input__4__ready),
    .input__4__valid(\input__4__valid$160 ),
    .input__5__payload(inputs__5__payload[4]),
    .input__5__ready(input__5__ready),
    .input__5__valid(\input__5__valid$162 ),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$319 ),
    .input__6__valid(\input__6__valid$164 ),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$328 ),
    .input__7__valid(\input__7__valid$166 ),
    .output__payload(\output__payload$171 ),
    .output__ready(\output__ready$172 ),
    .output__valid(\$signature__valid$168 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_1_arb  credit_counter_tx_east_vc_1_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(\input__0__ready$246 ),
    .input__0__valid(\input__0__valid$174 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(\input__1__ready$255 ),
    .input__1__valid(\input__1__valid$176 ),
    .input__2__payload(inputs__2__payload[4]),
    .input__2__ready(\input__2__ready$264 ),
    .input__2__valid(\input__2__valid$178 ),
    .input__3__payload(inputs__3__payload[4]),
    .input__3__ready(\input__3__ready$273 ),
    .input__3__valid(\input__3__valid$180 ),
    .input__4__payload(inputs__4__payload[4]),
    .input__4__ready(\input__4__ready$282 ),
    .input__4__valid(\input__4__valid$182 ),
    .input__5__payload(inputs__5__payload[4]),
    .input__5__ready(\input__5__ready$291 ),
    .input__5__valid(\input__5__valid$184 ),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$320 ),
    .input__6__valid(\input__6__valid$186 ),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$329 ),
    .input__7__valid(\input__7__valid$188 ),
    .output__payload(\output__payload$193 ),
    .output__ready(\output__ready$194 ),
    .output__valid(\$signature__valid$190 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_0_arb  credit_counter_tx_local_vc_0_arb (
    .clk(clk),
    .input__0__payload(inputs__2__payload[4]),
    .input__0__ready(\input__0__ready$259 ),
    .input__0__valid(input__0__valid),
    .input__1__payload(inputs__3__payload[4]),
    .input__1__ready(\input__1__ready$268 ),
    .input__1__valid(input__1__valid),
    .input__2__payload(inputs__4__payload[4]),
    .input__2__ready(\input__2__ready$277 ),
    .input__2__valid(input__2__valid),
    .input__3__payload(inputs__5__payload[4]),
    .input__3__ready(\input__3__ready$286 ),
    .input__3__valid(input__3__valid),
    .input__4__payload(inputs__6__payload[4]),
    .input__4__ready(\input__4__ready$295 ),
    .input__4__valid(input__4__valid),
    .input__5__payload(inputs__7__payload[4]),
    .input__5__ready(\input__5__ready$304 ),
    .input__5__valid(input__5__valid),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$313 ),
    .input__6__valid(input__6__valid),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$322 ),
    .input__7__valid(input__7__valid),
    .output__payload(output__payload),
    .output__ready(output__ready),
    .output__valid(\$signature__valid ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_1_arb  credit_counter_tx_local_vc_1_arb (
    .clk(clk),
    .input__0__payload(inputs__2__payload[4]),
    .input__0__ready(\input__0__ready$260 ),
    .input__0__valid(\input__0__valid$38 ),
    .input__1__payload(inputs__3__payload[4]),
    .input__1__ready(\input__1__ready$269 ),
    .input__1__valid(\input__1__valid$40 ),
    .input__2__payload(inputs__4__payload[4]),
    .input__2__ready(\input__2__ready$278 ),
    .input__2__valid(\input__2__valid$42 ),
    .input__3__payload(inputs__5__payload[4]),
    .input__3__ready(\input__3__ready$287 ),
    .input__3__valid(\input__3__valid$44 ),
    .input__4__payload(inputs__6__payload[4]),
    .input__4__ready(\input__4__ready$296 ),
    .input__4__valid(\input__4__valid$46 ),
    .input__5__payload(inputs__7__payload[4]),
    .input__5__ready(\input__5__ready$305 ),
    .input__5__valid(\input__5__valid$48 ),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$314 ),
    .input__6__valid(\input__6__valid$50 ),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$323 ),
    .input__7__valid(\input__7__valid$52 ),
    .output__payload(\output__payload$57 ),
    .output__ready(\output__ready$58 ),
    .output__valid(\$signature__valid$54 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:409" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north  credit_counter_tx_north (
    .clk(clk),
    .credit_in__payload(credit_in__payload),
    .credit_in__valid(credit_in__valid),
    .input__0__ready(\output__ready$84 ),
    .input__0__valid(\$signature__valid$80 ),
    .input__1__ready(\output__ready$106 ),
    .input__1__valid(\$signature__valid$102 ),
    .output__0__payload(\$signature__payload$82 ),
    .output__0__ready(output__0__ready),
    .output__0__valid(output__0__valid),
    .output__1__payload(\$signature__payload$104 ),
    .output__1__ready(output__1__ready),
    .output__1__valid(output__1__valid),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_0_arb  credit_counter_tx_north_vc_0_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(input__0__ready),
    .input__0__valid(\input__0__valid$60 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(input__1__ready),
    .input__1__valid(\input__1__valid$64 ),
    .input__2__payload(inputs__4__payload[4]),
    .input__2__ready(\input__2__ready$279 ),
    .input__2__valid(\input__2__valid$68 ),
    .input__3__payload(inputs__5__payload[4]),
    .input__3__ready(\input__3__ready$288 ),
    .input__3__valid(\input__3__valid$70 ),
    .input__4__payload(inputs__6__payload[4]),
    .input__4__ready(\input__4__ready$297 ),
    .input__4__valid(\input__4__valid$72 ),
    .input__5__payload(inputs__7__payload[4]),
    .input__5__ready(\input__5__ready$306 ),
    .input__5__valid(\input__5__valid$74 ),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$315 ),
    .input__6__valid(\input__6__valid$76 ),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$324 ),
    .input__7__valid(\input__7__valid$78 ),
    .output__payload(\output__payload$83 ),
    .output__ready(\output__ready$84 ),
    .output__valid(\$signature__valid$80 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_1_arb  credit_counter_tx_north_vc_1_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(\input__0__ready$242 ),
    .input__0__valid(\input__0__valid$86 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(\input__1__ready$251 ),
    .input__1__valid(\input__1__valid$88 ),
    .input__2__payload(inputs__4__payload[4]),
    .input__2__ready(\input__2__ready$280 ),
    .input__2__valid(\input__2__valid$90 ),
    .input__3__payload(inputs__5__payload[4]),
    .input__3__ready(\input__3__ready$289 ),
    .input__3__valid(\input__3__valid$92 ),
    .input__4__payload(inputs__6__payload[4]),
    .input__4__ready(\input__4__ready$298 ),
    .input__4__valid(\input__4__valid$94 ),
    .input__5__payload(inputs__7__payload[4]),
    .input__5__ready(\input__5__ready$307 ),
    .input__5__valid(\input__5__valid$96 ),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$316 ),
    .input__6__valid(\input__6__valid$98 ),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$325 ),
    .input__7__valid(\input__7__valid$100 ),
    .output__payload(\output__payload$105 ),
    .output__ready(\output__ready$106 ),
    .output__valid(\$signature__valid$102 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:409" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south  credit_counter_tx_south (
    .clk(clk),
    .credit_in__payload(\credit_in__payload$354 ),
    .credit_in__valid(\credit_in__valid$356 ),
    .input__0__ready(\output__ready$128 ),
    .input__0__valid(\$signature__valid$124 ),
    .input__1__ready(\output__ready$150 ),
    .input__1__valid(\$signature__valid$146 ),
    .output__0__payload(\$signature__payload$126 ),
    .output__0__ready(\output__0__ready$361 ),
    .output__0__valid(\output__0__valid$399 ),
    .output__1__payload(\$signature__payload$148 ),
    .output__1__ready(\output__1__ready$366 ),
    .output__1__valid(\output__1__valid$400 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_0_arb  credit_counter_tx_south_vc_0_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(\input__0__ready$243 ),
    .input__0__valid(\input__0__valid$108 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(\input__1__ready$252 ),
    .input__1__valid(\input__1__valid$110 ),
    .input__2__payload(inputs__2__payload[4]),
    .input__2__ready(input__2__ready),
    .input__2__valid(\input__2__valid$112 ),
    .input__3__payload(inputs__3__payload[4]),
    .input__3__ready(input__3__ready),
    .input__3__valid(\input__3__valid$114 ),
    .input__4__payload(inputs__6__payload[4]),
    .input__4__ready(\input__4__ready$299 ),
    .input__4__valid(\input__4__valid$116 ),
    .input__5__payload(inputs__7__payload[4]),
    .input__5__ready(\input__5__ready$308 ),
    .input__5__valid(\input__5__valid$118 ),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$317 ),
    .input__6__valid(\input__6__valid$120 ),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$326 ),
    .input__7__valid(\input__7__valid$122 ),
    .output__payload(\output__payload$127 ),
    .output__ready(\output__ready$128 ),
    .output__valid(\$signature__valid$124 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_1_arb  credit_counter_tx_south_vc_1_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(\input__0__ready$244 ),
    .input__0__valid(\input__0__valid$130 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(\input__1__ready$253 ),
    .input__1__valid(\input__1__valid$132 ),
    .input__2__payload(inputs__2__payload[4]),
    .input__2__ready(\input__2__ready$262 ),
    .input__2__valid(\input__2__valid$134 ),
    .input__3__payload(inputs__3__payload[4]),
    .input__3__ready(\input__3__ready$271 ),
    .input__3__valid(\input__3__valid$136 ),
    .input__4__payload(inputs__6__payload[4]),
    .input__4__ready(\input__4__ready$300 ),
    .input__4__valid(\input__4__valid$138 ),
    .input__5__payload(inputs__7__payload[4]),
    .input__5__ready(\input__5__ready$309 ),
    .input__5__valid(\input__5__valid$140 ),
    .input__6__payload(inputs__8__payload[4]),
    .input__6__ready(\input__6__ready$318 ),
    .input__6__valid(\input__6__valid$142 ),
    .input__7__payload(inputs__9__payload[4]),
    .input__7__ready(\input__7__ready$327 ),
    .input__7__valid(\input__7__valid$144 ),
    .output__payload(\output__payload$149 ),
    .output__ready(\output__ready$150 ),
    .output__valid(\$signature__valid$146 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:409" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west  credit_counter_tx_west (
    .clk(clk),
    .credit_in__payload(\credit_in__payload$382 ),
    .credit_in__valid(\credit_in__valid$384 ),
    .input__0__ready(\output__ready$216 ),
    .input__0__valid(\$signature__valid$212 ),
    .input__1__ready(\output__ready$238 ),
    .input__1__valid(\$signature__valid$234 ),
    .output__0__ready(\output__0__ready$389 ),
    .output__0__valid(\output__0__valid$403 ),
    .output__1__ready(\output__1__ready$394 ),
    .output__1__valid(\output__1__valid$404 ),
    .\port$216$0 (\$73 ),
    .\port$234$0 (\$82 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_0_arb  credit_counter_tx_west_vc_0_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(\input__0__ready$247 ),
    .input__0__valid(\input__0__valid$196 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(\input__1__ready$256 ),
    .input__1__valid(\input__1__valid$198 ),
    .input__2__payload(inputs__2__payload[4]),
    .input__2__ready(\input__2__ready$265 ),
    .input__2__valid(\input__2__valid$200 ),
    .input__3__payload(inputs__3__payload[4]),
    .input__3__ready(\input__3__ready$274 ),
    .input__3__valid(\input__3__valid$202 ),
    .input__4__payload(inputs__4__payload[4]),
    .input__4__ready(\input__4__ready$283 ),
    .input__4__valid(\input__4__valid$204 ),
    .input__5__payload(inputs__5__payload[4]),
    .input__5__ready(\input__5__ready$292 ),
    .input__5__valid(\input__5__valid$206 ),
    .input__6__payload(inputs__6__payload[4]),
    .input__6__ready(input__6__ready),
    .input__6__valid(\input__6__valid$208 ),
    .input__7__payload(inputs__7__payload[4]),
    .input__7__ready(input__7__ready),
    .input__7__valid(\input__7__valid$210 ),
    .output__payload(\output__payload$215 ),
    .output__ready(\output__ready$216 ),
    .output__valid(\$signature__valid$212 ),
    .rst(rst)
  );
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/memory_mapped_router.py:384" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_1_arb  credit_counter_tx_west_vc_1_arb (
    .clk(clk),
    .input__0__payload(inputs__0__payload[4]),
    .input__0__ready(\input__0__ready$248 ),
    .input__0__valid(\input__0__valid$218 ),
    .input__1__payload(inputs__1__payload[4]),
    .input__1__ready(\input__1__ready$257 ),
    .input__1__valid(\input__1__valid$220 ),
    .input__2__payload(inputs__2__payload[4]),
    .input__2__ready(\input__2__ready$266 ),
    .input__2__valid(\input__2__valid$222 ),
    .input__3__payload(inputs__3__payload[4]),
    .input__3__ready(\input__3__ready$275 ),
    .input__3__valid(\input__3__valid$224 ),
    .input__4__payload(inputs__4__payload[4]),
    .input__4__ready(\input__4__ready$284 ),
    .input__4__valid(\input__4__valid$226 ),
    .input__5__payload(inputs__5__payload[4]),
    .input__5__ready(\input__5__ready$293 ),
    .input__5__valid(\input__5__valid$228 ),
    .input__6__payload(inputs__6__payload[4]),
    .input__6__ready(\input__6__ready$302 ),
    .input__6__valid(\input__6__valid$230 ),
    .input__7__payload(inputs__7__payload[4]),
    .input__7__ready(\input__7__ready$311 ),
    .input__7__valid(\input__7__valid$232 ),
    .output__payload(\output__payload$237 ),
    .output__ready(\output__ready$238 ),
    .output__valid(\$signature__valid$234 ),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (output__payload[3:1])
      3'h0:
          \$signature__payload  = 4'h2;
      3'h1:
          \$signature__payload  = 4'h3;
      3'h2:
          \$signature__payload  = 4'h4;
      3'h3:
          \$signature__payload  = 4'h5;
      3'h4:
          \$signature__payload  = 4'h6;
      3'h5:
          \$signature__payload  = 4'h7;
      3'h6:
          \$signature__payload  = 4'h8;
      3'h7:
          \$signature__payload  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$57 [3:1])
      3'h0:
          \$signature__payload$56  = 4'h2;
      3'h1:
          \$signature__payload$56  = 4'h3;
      3'h2:
          \$signature__payload$56  = 4'h4;
      3'h3:
          \$signature__payload$56  = 4'h5;
      3'h4:
          \$signature__payload$56  = 4'h6;
      3'h5:
          \$signature__payload$56  = 4'h7;
      3'h6:
          \$signature__payload$56  = 4'h8;
      3'h7:
          \$signature__payload$56  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$83 [3:1])
      3'h0:
          \$signature__payload$82  = 4'h0;
      3'h1:
          \$signature__payload$82  = 4'h1;
      3'h2:
          \$signature__payload$82  = 4'h4;
      3'h3:
          \$signature__payload$82  = 4'h5;
      3'h4:
          \$signature__payload$82  = 4'h6;
      3'h5:
          \$signature__payload$82  = 4'h7;
      3'h6:
          \$signature__payload$82  = 4'h8;
      3'h7:
          \$signature__payload$82  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$105 [3:1])
      3'h0:
          \$signature__payload$104  = 4'h0;
      3'h1:
          \$signature__payload$104  = 4'h1;
      3'h2:
          \$signature__payload$104  = 4'h4;
      3'h3:
          \$signature__payload$104  = 4'h5;
      3'h4:
          \$signature__payload$104  = 4'h6;
      3'h5:
          \$signature__payload$104  = 4'h7;
      3'h6:
          \$signature__payload$104  = 4'h8;
      3'h7:
          \$signature__payload$104  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$127 [3:1])
      3'h0:
          \$signature__payload$126  = 4'h0;
      3'h1:
          \$signature__payload$126  = 4'h1;
      3'h2:
          \$signature__payload$126  = 4'h2;
      3'h3:
          \$signature__payload$126  = 4'h3;
      3'h4:
          \$signature__payload$126  = 4'h6;
      3'h5:
          \$signature__payload$126  = 4'h7;
      3'h6:
          \$signature__payload$126  = 4'h8;
      3'h7:
          \$signature__payload$126  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$149 [3:1])
      3'h0:
          \$signature__payload$148  = 4'h0;
      3'h1:
          \$signature__payload$148  = 4'h1;
      3'h2:
          \$signature__payload$148  = 4'h2;
      3'h3:
          \$signature__payload$148  = 4'h3;
      3'h4:
          \$signature__payload$148  = 4'h6;
      3'h5:
          \$signature__payload$148  = 4'h7;
      3'h6:
          \$signature__payload$148  = 4'h8;
      3'h7:
          \$signature__payload$148  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$171 [3:1])
      3'h0:
          \$signature__payload$170  = 4'h0;
      3'h1:
          \$signature__payload$170  = 4'h1;
      3'h2:
          \$signature__payload$170  = 4'h2;
      3'h3:
          \$signature__payload$170  = 4'h3;
      3'h4:
          \$signature__payload$170  = 4'h4;
      3'h5:
          \$signature__payload$170  = 4'h5;
      3'h6:
          \$signature__payload$170  = 4'h8;
      3'h7:
          \$signature__payload$170  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$193 [3:1])
      3'h0:
          \$signature__payload$192  = 4'h0;
      3'h1:
          \$signature__payload$192  = 4'h1;
      3'h2:
          \$signature__payload$192  = 4'h2;
      3'h3:
          \$signature__payload$192  = 4'h3;
      3'h4:
          \$signature__payload$192  = 4'h4;
      3'h5:
          \$signature__payload$192  = 4'h5;
      3'h6:
          \$signature__payload$192  = 4'h8;
      3'h7:
          \$signature__payload$192  = 4'h9;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$215 [3:1])
      3'h0:
          \$73  = 3'h0;
      3'h1:
          \$73  = 3'h1;
      3'h2:
          \$73  = 3'h2;
      3'h3:
          \$73  = 3'h3;
      3'h4:
          \$73  = 3'h4;
      3'h5:
          \$73  = 3'h5;
      3'h6:
          \$73  = 3'h6;
      3'h7:
          \$73  = 3'h7;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez (\output__payload$237 [3:1])
      3'h0:
          \$82  = 3'h0;
      3'h1:
          \$82  = 3'h1;
      3'h2:
          \$82  = 3'h2;
      3'h3:
          \$82  = 3'h3;
      3'h4:
          \$82  = 3'h4;
      3'h5:
          \$82  = 3'h5;
      3'h6:
          \$82  = 3'h6;
      3'h7:
          \$82  = 3'h7;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    output__ready = 1'h0;
    casez (\$signature__payload )
      4'h0:
          output__ready = outputs__0__ready;
      4'h1:
          output__ready = outputs__1__ready;
      4'h2:
          output__ready = outputs__2__ready;
      4'h3:
          output__ready = outputs__3__ready;
      4'h4:
          output__ready = outputs__4__ready;
      4'h5:
          output__ready = outputs__5__ready;
      4'h6:
          output__ready = outputs__6__ready;
      4'h7:
          output__ready = outputs__7__ready;
      4'h8:
          output__ready = outputs__8__ready;
      4'h9:
          output__ready = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    \output__ready$58  = 1'h0;
    casez (\$signature__payload$56 )
      4'h0:
          \output__ready$58  = outputs__0__ready;
      4'h1:
          \output__ready$58  = outputs__1__ready;
      4'h2:
          \output__ready$58  = outputs__2__ready;
      4'h3:
          \output__ready$58  = outputs__3__ready;
      4'h4:
          \output__ready$58  = outputs__4__ready;
      4'h5:
          \output__ready$58  = outputs__5__ready;
      4'h6:
          \output__ready$58  = outputs__6__ready;
      4'h7:
          \output__ready$58  = outputs__7__ready;
      4'h8:
          \output__ready$58  = outputs__8__ready;
      4'h9:
          \output__ready$58  = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    output__0__ready = 1'h0;
    casez (\$signature__payload$82 )
      4'h0:
          output__0__ready = outputs__0__ready;
      4'h1:
          output__0__ready = outputs__1__ready;
      4'h2:
          output__0__ready = outputs__2__ready;
      4'h3:
          output__0__ready = outputs__3__ready;
      4'h4:
          output__0__ready = outputs__4__ready;
      4'h5:
          output__0__ready = outputs__5__ready;
      4'h6:
          output__0__ready = outputs__6__ready;
      4'h7:
          output__0__ready = outputs__7__ready;
      4'h8:
          output__0__ready = outputs__8__ready;
      4'h9:
          output__0__ready = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    output__1__ready = 1'h0;
    casez (\$signature__payload$104 )
      4'h0:
          output__1__ready = outputs__0__ready;
      4'h1:
          output__1__ready = outputs__1__ready;
      4'h2:
          output__1__ready = outputs__2__ready;
      4'h3:
          output__1__ready = outputs__3__ready;
      4'h4:
          output__1__ready = outputs__4__ready;
      4'h5:
          output__1__ready = outputs__5__ready;
      4'h6:
          output__1__ready = outputs__6__ready;
      4'h7:
          output__1__ready = outputs__7__ready;
      4'h8:
          output__1__ready = outputs__8__ready;
      4'h9:
          output__1__ready = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    \output__0__ready$361  = 1'h0;
    casez (\$signature__payload$126 )
      4'h0:
          \output__0__ready$361  = outputs__0__ready;
      4'h1:
          \output__0__ready$361  = outputs__1__ready;
      4'h2:
          \output__0__ready$361  = outputs__2__ready;
      4'h3:
          \output__0__ready$361  = outputs__3__ready;
      4'h4:
          \output__0__ready$361  = outputs__4__ready;
      4'h5:
          \output__0__ready$361  = outputs__5__ready;
      4'h6:
          \output__0__ready$361  = outputs__6__ready;
      4'h7:
          \output__0__ready$361  = outputs__7__ready;
      4'h8:
          \output__0__ready$361  = outputs__8__ready;
      4'h9:
          \output__0__ready$361  = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    \output__1__ready$366  = 1'h0;
    casez (\$signature__payload$148 )
      4'h0:
          \output__1__ready$366  = outputs__0__ready;
      4'h1:
          \output__1__ready$366  = outputs__1__ready;
      4'h2:
          \output__1__ready$366  = outputs__2__ready;
      4'h3:
          \output__1__ready$366  = outputs__3__ready;
      4'h4:
          \output__1__ready$366  = outputs__4__ready;
      4'h5:
          \output__1__ready$366  = outputs__5__ready;
      4'h6:
          \output__1__ready$366  = outputs__6__ready;
      4'h7:
          \output__1__ready$366  = outputs__7__ready;
      4'h8:
          \output__1__ready$366  = outputs__8__ready;
      4'h9:
          \output__1__ready$366  = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    \output__0__ready$375  = 1'h0;
    casez (\$signature__payload$170 )
      4'h0:
          \output__0__ready$375  = outputs__0__ready;
      4'h1:
          \output__0__ready$375  = outputs__1__ready;
      4'h2:
          \output__0__ready$375  = outputs__2__ready;
      4'h3:
          \output__0__ready$375  = outputs__3__ready;
      4'h4:
          \output__0__ready$375  = outputs__4__ready;
      4'h5:
          \output__0__ready$375  = outputs__5__ready;
      4'h6:
          \output__0__ready$375  = outputs__6__ready;
      4'h7:
          \output__0__ready$375  = outputs__7__ready;
      4'h8:
          \output__0__ready$375  = outputs__8__ready;
      4'h9:
          \output__0__ready$375  = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    \output__1__ready$380  = 1'h0;
    casez (\$signature__payload$192 )
      4'h0:
          \output__1__ready$380  = outputs__0__ready;
      4'h1:
          \output__1__ready$380  = outputs__1__ready;
      4'h2:
          \output__1__ready$380  = outputs__2__ready;
      4'h3:
          \output__1__ready$380  = outputs__3__ready;
      4'h4:
          \output__1__ready$380  = outputs__4__ready;
      4'h5:
          \output__1__ready$380  = outputs__5__ready;
      4'h6:
          \output__1__ready$380  = outputs__6__ready;
      4'h7:
          \output__1__ready$380  = outputs__7__ready;
      4'h8:
          \output__1__ready$380  = outputs__8__ready;
      4'h9:
          \output__1__ready$380  = outputs__9__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez ({ 1'h0, \$73  })
      4'h0:
          \output__0__ready$389  = outputs__0__ready;
      4'h1:
          \output__0__ready$389  = outputs__1__ready;
      4'h2:
          \output__0__ready$389  = outputs__2__ready;
      4'h3:
          \output__0__ready$389  = outputs__3__ready;
      4'h4:
          \output__0__ready$389  = outputs__4__ready;
      4'h5:
          \output__0__ready$389  = outputs__5__ready;
      4'h6:
          \output__0__ready$389  = outputs__6__ready;
      4'h7:
          \output__0__ready$389  = outputs__7__ready;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$33 ) begin end
    (* full_case = 32'd1 *)
    casez ({ 1'h0, \$82  })
      4'h0:
          \output__1__ready$394  = outputs__0__ready;
      4'h1:
          \output__1__ready$394  = outputs__1__ready;
      4'h2:
          \output__1__ready$394  = outputs__2__ready;
      4'h3:
          \output__1__ready$394  = outputs__3__ready;
      4'h4:
          \output__1__ready$394  = outputs__4__ready;
      4'h5:
          \output__1__ready$394  = outputs__5__ready;
      4'h6:
          \output__1__ready$394  = outputs__6__ready;
      4'h7:
          \output__1__ready$394  = outputs__7__ready;
    endcase
  end
  assign input__0__payload = inputs__2__payload[4];
  assign input__1__payload = inputs__3__payload[4];
  assign input__2__payload = inputs__4__payload[4];
  assign input__3__payload = inputs__5__payload[4];
  assign input__4__payload = inputs__6__payload[4];
  assign input__5__payload = inputs__7__payload[4];
  assign input__6__payload = inputs__8__payload[4];
  assign input__7__payload = inputs__9__payload[4];
  assign output__valid = \$signature__valid ;
  assign \$signature__ready  = output__ready;
  assign \input__0__payload$39  = inputs__2__payload[4];
  assign \input__1__payload$41  = inputs__3__payload[4];
  assign \input__2__payload$43  = inputs__4__payload[4];
  assign \input__3__payload$45  = inputs__5__payload[4];
  assign \input__4__payload$47  = inputs__6__payload[4];
  assign \input__5__payload$49  = inputs__7__payload[4];
  assign \input__6__payload$51  = inputs__8__payload[4];
  assign \input__7__payload$53  = inputs__9__payload[4];
  assign \output__valid$55  = \$signature__valid$54 ;
  assign \$signature__ready$59  = \output__ready$58 ;
  assign \input__0__payload$63  = inputs__0__payload[4];
  assign \input__1__payload$67  = inputs__1__payload[4];
  assign \input__2__payload$69  = inputs__4__payload[4];
  assign \input__3__payload$71  = inputs__5__payload[4];
  assign \input__4__payload$73  = inputs__6__payload[4];
  assign \input__5__payload$75  = inputs__7__payload[4];
  assign \input__6__payload$77  = inputs__8__payload[4];
  assign \input__7__payload$79  = inputs__9__payload[4];
  assign \output__valid$81  = \$signature__valid$80 ;
  assign \$signature__ready$85  = \output__ready$84 ;
  assign \input__0__payload$87  = inputs__0__payload[4];
  assign \input__1__payload$89  = inputs__1__payload[4];
  assign \input__2__payload$91  = inputs__4__payload[4];
  assign \input__3__payload$93  = inputs__5__payload[4];
  assign \input__4__payload$95  = inputs__6__payload[4];
  assign \input__5__payload$97  = inputs__7__payload[4];
  assign \input__6__payload$99  = inputs__8__payload[4];
  assign \input__7__payload$101  = inputs__9__payload[4];
  assign \output__valid$103  = \$signature__valid$102 ;
  assign \$signature__ready$107  = \output__ready$106 ;
  assign \input__0__payload$109  = inputs__0__payload[4];
  assign \input__1__payload$111  = inputs__1__payload[4];
  assign \input__2__payload$113  = inputs__2__payload[4];
  assign \input__3__payload$115  = inputs__3__payload[4];
  assign \input__4__payload$117  = inputs__6__payload[4];
  assign \input__5__payload$119  = inputs__7__payload[4];
  assign \input__6__payload$121  = inputs__8__payload[4];
  assign \input__7__payload$123  = inputs__9__payload[4];
  assign \output__valid$125  = \$signature__valid$124 ;
  assign \$signature__ready$129  = \output__ready$128 ;
  assign \input__0__payload$131  = inputs__0__payload[4];
  assign \input__1__payload$133  = inputs__1__payload[4];
  assign \input__2__payload$135  = inputs__2__payload[4];
  assign \input__3__payload$137  = inputs__3__payload[4];
  assign \input__4__payload$139  = inputs__6__payload[4];
  assign \input__5__payload$141  = inputs__7__payload[4];
  assign \input__6__payload$143  = inputs__8__payload[4];
  assign \input__7__payload$145  = inputs__9__payload[4];
  assign \output__valid$147  = \$signature__valid$146 ;
  assign \$signature__ready$151  = \output__ready$150 ;
  assign \input__0__payload$153  = inputs__0__payload[4];
  assign \input__1__payload$155  = inputs__1__payload[4];
  assign \input__2__payload$157  = inputs__2__payload[4];
  assign \input__3__payload$159  = inputs__3__payload[4];
  assign \input__4__payload$161  = inputs__4__payload[4];
  assign \input__5__payload$163  = inputs__5__payload[4];
  assign \input__6__payload$165  = inputs__8__payload[4];
  assign \input__7__payload$167  = inputs__9__payload[4];
  assign \output__valid$169  = \$signature__valid$168 ;
  assign \$signature__ready$173  = \output__ready$172 ;
  assign \input__0__payload$175  = inputs__0__payload[4];
  assign \input__1__payload$177  = inputs__1__payload[4];
  assign \input__2__payload$179  = inputs__2__payload[4];
  assign \input__3__payload$181  = inputs__3__payload[4];
  assign \input__4__payload$183  = inputs__4__payload[4];
  assign \input__5__payload$185  = inputs__5__payload[4];
  assign \input__6__payload$187  = inputs__8__payload[4];
  assign \input__7__payload$189  = inputs__9__payload[4];
  assign \output__valid$191  = \$signature__valid$190 ;
  assign \$signature__ready$195  = \output__ready$194 ;
  assign \input__0__payload$197  = inputs__0__payload[4];
  assign \input__1__payload$199  = inputs__1__payload[4];
  assign \input__2__payload$201  = inputs__2__payload[4];
  assign \input__3__payload$203  = inputs__3__payload[4];
  assign \input__4__payload$205  = inputs__4__payload[4];
  assign \input__5__payload$207  = inputs__5__payload[4];
  assign \input__6__payload$209  = inputs__6__payload[4];
  assign \input__7__payload$211  = inputs__7__payload[4];
  assign \output__valid$213  = \$signature__valid$212 ;
  assign \$signature__payload$214  = { 1'h0, \$73  };
  assign \$signature__ready$217  = \output__ready$216 ;
  assign \input__0__payload$219  = inputs__0__payload[4];
  assign \input__1__payload$221  = inputs__1__payload[4];
  assign \input__2__payload$223  = inputs__2__payload[4];
  assign \input__3__payload$225  = inputs__3__payload[4];
  assign \input__4__payload$227  = inputs__4__payload[4];
  assign \input__5__payload$229  = inputs__5__payload[4];
  assign \input__6__payload$231  = inputs__6__payload[4];
  assign \input__7__payload$233  = inputs__7__payload[4];
  assign \output__valid$235  = \$signature__valid$234 ;
  assign \$signature__payload$236  = { 1'h0, \$82  };
  assign \$signature__ready$239  = \output__ready$238 ;
  assign credit__0__payload = credit_in__payload;
  assign credit__0__valid = credit_in__valid;
  assign \input__0__payload$344  = \$signature__payload$82 ;
  assign \input__0__ready$345  = \output__ready$84 ;
  assign \input__0__valid$346  = \$signature__valid$80 ;
  assign output__0__payload = \$signature__payload$82 ;
  assign \input__1__payload$349  = \$signature__payload$104 ;
  assign \input__1__ready$350  = \output__ready$106 ;
  assign \input__1__valid$351  = \$signature__valid$102 ;
  assign output__1__payload = \$signature__payload$104 ;
  assign credit__1__payload = \credit_in__payload$354 ;
  assign credit__1__valid = \credit_in__valid$356 ;
  assign \input__0__payload$358  = \$signature__payload$126 ;
  assign \input__0__ready$359  = \output__ready$128 ;
  assign \input__0__valid$360  = \$signature__valid$124 ;
  assign \output__0__payload$362  = \$signature__payload$126 ;
  assign \input__1__payload$363  = \$signature__payload$148 ;
  assign \input__1__ready$364  = \output__ready$150 ;
  assign \input__1__valid$365  = \$signature__valid$146 ;
  assign \output__1__payload$367  = \$signature__payload$148 ;
  assign credit__2__payload = \credit_in__payload$368 ;
  assign credit__2__valid = \credit_in__valid$370 ;
  assign \input__0__payload$372  = \$signature__payload$170 ;
  assign \input__0__ready$373  = \output__ready$172 ;
  assign \input__0__valid$374  = \$signature__valid$168 ;
  assign \output__0__payload$376  = \$signature__payload$170 ;
  assign \input__1__payload$377  = \$signature__payload$192 ;
  assign \input__1__ready$378  = \output__ready$194 ;
  assign \input__1__valid$379  = \$signature__valid$190 ;
  assign \output__1__payload$381  = \$signature__payload$192 ;
  assign credit__3__payload = \credit_in__payload$382 ;
  assign credit__3__valid = \credit_in__valid$384 ;
  assign \input__0__payload$386  = { 1'h0, \$73  };
  assign \input__0__ready$387  = \output__ready$216 ;
  assign \input__0__valid$388  = \$signature__valid$212 ;
  assign \output__0__payload$390  = { 1'h0, \$73  };
  assign \input__1__payload$391  = { 1'h0, \$82  };
  assign \input__1__ready$392  = \output__ready$238 ;
  assign \input__1__valid$393  = \$signature__valid$234 ;
  assign \output__1__payload$395  = { 1'h0, \$82  };
  assign \inputs__2__payload.target  = inputs__2__payload[3:0];
  assign \inputs__2__payload.target.port  = inputs__2__payload[2:0];
  assign \inputs__2__payload.target.vc_id  = inputs__2__payload[3];
  assign \inputs__2__payload.last  = inputs__2__payload[4];
  assign \inputs__3__payload.target  = inputs__3__payload[3:0];
  assign \inputs__3__payload.target.port  = inputs__3__payload[2:0];
  assign \inputs__3__payload.target.vc_id  = inputs__3__payload[3];
  assign \inputs__3__payload.last  = inputs__3__payload[4];
  assign \inputs__4__payload.target  = inputs__4__payload[3:0];
  assign \inputs__4__payload.target.port  = inputs__4__payload[2:0];
  assign \inputs__4__payload.target.vc_id  = inputs__4__payload[3];
  assign \inputs__4__payload.last  = inputs__4__payload[4];
  assign \inputs__5__payload.target  = inputs__5__payload[3:0];
  assign \inputs__5__payload.target.port  = inputs__5__payload[2:0];
  assign \inputs__5__payload.target.vc_id  = inputs__5__payload[3];
  assign \inputs__5__payload.last  = inputs__5__payload[4];
  assign \inputs__6__payload.target  = inputs__6__payload[3:0];
  assign \inputs__6__payload.target.port  = inputs__6__payload[2:0];
  assign \inputs__6__payload.target.vc_id  = inputs__6__payload[3];
  assign \inputs__6__payload.last  = inputs__6__payload[4];
  assign \inputs__7__payload.target  = inputs__7__payload[3:0];
  assign \inputs__7__payload.target.port  = inputs__7__payload[2:0];
  assign \inputs__7__payload.target.vc_id  = inputs__7__payload[3];
  assign \inputs__7__payload.last  = inputs__7__payload[4];
  assign \inputs__8__payload.target  = inputs__8__payload[3:0];
  assign \inputs__8__payload.target.port  = inputs__8__payload[2:0];
  assign \inputs__8__payload.target.vc_id  = inputs__8__payload[3];
  assign \inputs__8__payload.last  = inputs__8__payload[4];
  assign \inputs__9__payload.target  = inputs__9__payload[3:0];
  assign \inputs__9__payload.target.port  = inputs__9__payload[2:0];
  assign \inputs__9__payload.target.vc_id  = inputs__9__payload[3];
  assign \inputs__9__payload.last  = inputs__9__payload[4];
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign \output__payload$57.last  = \output__payload$57 [0];
  assign \output__payload$57.src  = \output__payload$57 [3:1];
  assign \inputs__0__payload.target  = inputs__0__payload[3:0];
  assign \inputs__0__payload.target.port  = inputs__0__payload[2:0];
  assign \inputs__0__payload.target.vc_id  = inputs__0__payload[3];
  assign \inputs__0__payload.last  = inputs__0__payload[4];
  assign \inputs__1__payload.target  = inputs__1__payload[3:0];
  assign \inputs__1__payload.target.port  = inputs__1__payload[2:0];
  assign \inputs__1__payload.target.vc_id  = inputs__1__payload[3];
  assign \inputs__1__payload.last  = inputs__1__payload[4];
  assign \output__payload$83.last  = \output__payload$83 [0];
  assign \output__payload$83.src  = \output__payload$83 [3:1];
  assign \output__payload$105.last  = \output__payload$105 [0];
  assign \output__payload$105.src  = \output__payload$105 [3:1];
  assign \output__payload$127.last  = \output__payload$127 [0];
  assign \output__payload$127.src  = \output__payload$127 [3:1];
  assign \output__payload$149.last  = \output__payload$149 [0];
  assign \output__payload$149.src  = \output__payload$149 [3:1];
  assign \output__payload$171.last  = \output__payload$171 [0];
  assign \output__payload$171.src  = \output__payload$171 [3:1];
  assign \output__payload$193.last  = \output__payload$193 [0];
  assign \output__payload$193.src  = \output__payload$193 [3:1];
  assign \output__payload$215.last  = \output__payload$215 [0];
  assign \output__payload$215.src  = \output__payload$215 [3:1];
  assign \output__payload$237.last  = \output__payload$237 [0];
  assign \output__payload$237.src  = \output__payload$237 [3:1];
  assign \credit_in__payload[0]  = credit_in__payload[5:0];
  assign \credit_in__payload[1]  = credit_in__payload[11:6];
  assign \credit__0__payload[0]  = credit_in__payload[5:0];
  assign \credit__0__payload[1]  = credit_in__payload[11:6];
  assign \credit_in__payload$354[0]  = \credit_in__payload$354 [5:0];
  assign \credit_in__payload$354[1]  = \credit_in__payload$354 [11:6];
  assign \credit__1__payload[0]  = \credit_in__payload$354 [5:0];
  assign \credit__1__payload[1]  = \credit_in__payload$354 [11:6];
  assign \credit_in__payload$368[0]  = \credit_in__payload$368 [5:0];
  assign \credit_in__payload$368[1]  = \credit_in__payload$368 [11:6];
  assign \credit__2__payload[0]  = \credit_in__payload$368 [5:0];
  assign \credit__2__payload[1]  = \credit_in__payload$368 [11:6];
  assign \credit_in__payload$382[0]  = \credit_in__payload$382 [5:0];
  assign \credit_in__payload$382[1]  = \credit_in__payload$382 [11:6];
  assign \credit__3__payload[0]  = \credit_in__payload$382 [5:0];
  assign \credit__3__payload[1]  = \credit_in__payload$382 [11:6];
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:832" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east (credit_in__valid, clk, rst, output__0__payload, output__1__payload, output__0__ready, output__1__ready, output__0__valid, input__0__ready, output__1__valid, input__1__ready, input__0__valid, input__1__valid, credit_in__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$34  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  reg [5:0] \$22 ;
  reg [5:0] \$23 ;
  reg [5:0] \$24 ;
  reg [5:0] \$25 ;
  wire [6:0] \$3 ;
  wire \$4 ;
  wire [6:0] \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  input [11:0] credit_in__payload;
  wire [11:0] credit_in__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit_in__valid;
  wire credit_in__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input [3:0] output__0__payload;
  wire [3:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input [3:0] output__1__payload;
  wire [3:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_1 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_1 = 6'h00;
  assign \$2  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__0__ready;
  assign \$3  = write_ptr_0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$4  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__1__ready;
  assign \$5  = write_ptr_1 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$6  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$7  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$8  = \$6  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$7 ;
  assign \$9  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$8 ;
  assign output__0__valid = input__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$9 ;
  assign \$10  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$11  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$12  = \$10  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$11 ;
  assign \$13  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$12 ;
  assign input__0__ready = output__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$13 ;
  assign \$14  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$15  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$16  = \$14  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$15 ;
  assign \$17  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$16 ;
  assign output__1__valid = input__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$17 ;
  assign \$18  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$19  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$20  = \$18  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$19 ;
  assign \$21  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$20 ;
  assign input__1__ready = output__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$21 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_0 <= \$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_1 <= \$23 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_0 <= \$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_1 <= \$25 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$34 ) begin end
    \$22  = read_ptr_0;
    if (\$1 ) begin
      \$22  = credit_in__payload[5:0];
    end
    if (rst) begin
      \$22  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$34 ) begin end
    \$23  = read_ptr_1;
    if (\$1 ) begin
      \$23  = credit_in__payload[11:6];
    end
    if (rst) begin
      \$23  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$34 ) begin end
    \$24  = write_ptr_0;
    if (\$2 ) begin
      \$24  = \$3 [5:0];
    end
    if (rst) begin
      \$24  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$34 ) begin end
    \$25  = write_ptr_1;
    if (\$4 ) begin
      \$25  = \$5 [5:0];
    end
    if (rst) begin
      \$25  = 6'h00;
    end
  end
  assign input__0__payload = output__0__payload;
  assign input__1__payload = output__1__payload;
  assign \credit_in__payload[0]  = credit_in__payload[5:0];
  assign \credit_in__payload[1]  = credit_in__payload[11:6];
  assign \$1  = credit_in__valid;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_0_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$35  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_0_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$35 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_0_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$36  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$36 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$36 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_1_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$37  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_1_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$37 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_east_vc_1_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$38  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$38 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$38 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_0_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$39  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_0_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$39 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_0_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$40  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$40 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$40 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_1_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$41  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_1_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$41 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_local_vc_1_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$42  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$42 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$42 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:832" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north (credit_in__valid, clk, rst, output__0__payload, output__1__payload, output__0__ready, output__1__ready, output__0__valid, input__0__ready, output__1__valid, input__1__ready, input__0__valid, input__1__valid, credit_in__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$43  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  reg [5:0] \$22 ;
  reg [5:0] \$23 ;
  reg [5:0] \$24 ;
  reg [5:0] \$25 ;
  wire [6:0] \$3 ;
  wire \$4 ;
  wire [6:0] \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  input [11:0] credit_in__payload;
  wire [11:0] credit_in__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit_in__valid;
  wire credit_in__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input [3:0] output__0__payload;
  wire [3:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input [3:0] output__1__payload;
  wire [3:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_1 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_1 = 6'h00;
  assign \$2  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__0__ready;
  assign \$3  = write_ptr_0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$4  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__1__ready;
  assign \$5  = write_ptr_1 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$6  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$7  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$8  = \$6  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$7 ;
  assign \$9  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$8 ;
  assign output__0__valid = input__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$9 ;
  assign \$10  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$11  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$12  = \$10  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$11 ;
  assign \$13  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$12 ;
  assign input__0__ready = output__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$13 ;
  assign \$14  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$15  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$16  = \$14  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$15 ;
  assign \$17  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$16 ;
  assign output__1__valid = input__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$17 ;
  assign \$18  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$19  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$20  = \$18  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$19 ;
  assign \$21  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$20 ;
  assign input__1__ready = output__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$21 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_0 <= \$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_1 <= \$23 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_0 <= \$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_1 <= \$25 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$43 ) begin end
    \$22  = read_ptr_0;
    if (\$1 ) begin
      \$22  = credit_in__payload[5:0];
    end
    if (rst) begin
      \$22  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$43 ) begin end
    \$23  = read_ptr_1;
    if (\$1 ) begin
      \$23  = credit_in__payload[11:6];
    end
    if (rst) begin
      \$23  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$43 ) begin end
    \$24  = write_ptr_0;
    if (\$2 ) begin
      \$24  = \$3 [5:0];
    end
    if (rst) begin
      \$24  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$43 ) begin end
    \$25  = write_ptr_1;
    if (\$4 ) begin
      \$25  = \$5 [5:0];
    end
    if (rst) begin
      \$25  = 6'h00;
    end
  end
  assign input__0__payload = output__0__payload;
  assign input__1__payload = output__1__payload;
  assign \credit_in__payload[0]  = credit_in__payload[5:0];
  assign \credit_in__payload[1]  = credit_in__payload[11:6];
  assign \$1  = credit_in__valid;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_0_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$44  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_0_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$44 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_0_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$45  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$45 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$45 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_1_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$46  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_1_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$46 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_north_vc_1_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$47  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$47 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$47 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:832" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south (credit_in__valid, clk, rst, output__0__payload, output__1__payload, output__0__ready, output__1__ready, output__0__valid, input__0__ready, output__1__valid, input__1__ready, input__0__valid, input__1__valid, credit_in__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$48  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  reg [5:0] \$22 ;
  reg [5:0] \$23 ;
  reg [5:0] \$24 ;
  reg [5:0] \$25 ;
  wire [6:0] \$3 ;
  wire \$4 ;
  wire [6:0] \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  input [11:0] credit_in__payload;
  wire [11:0] credit_in__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit_in__valid;
  wire credit_in__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input [3:0] output__0__payload;
  wire [3:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input [3:0] output__1__payload;
  wire [3:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_1 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_1 = 6'h00;
  assign \$2  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__0__ready;
  assign \$3  = write_ptr_0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$4  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__1__ready;
  assign \$5  = write_ptr_1 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$6  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$7  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$8  = \$6  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$7 ;
  assign \$9  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$8 ;
  assign output__0__valid = input__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$9 ;
  assign \$10  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$11  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$12  = \$10  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$11 ;
  assign \$13  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$12 ;
  assign input__0__ready = output__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$13 ;
  assign \$14  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$15  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$16  = \$14  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$15 ;
  assign \$17  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$16 ;
  assign output__1__valid = input__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$17 ;
  assign \$18  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$19  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$20  = \$18  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$19 ;
  assign \$21  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$20 ;
  assign input__1__ready = output__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$21 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_0 <= \$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_1 <= \$23 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_0 <= \$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_1 <= \$25 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$48 ) begin end
    \$22  = read_ptr_0;
    if (\$1 ) begin
      \$22  = credit_in__payload[5:0];
    end
    if (rst) begin
      \$22  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$48 ) begin end
    \$23  = read_ptr_1;
    if (\$1 ) begin
      \$23  = credit_in__payload[11:6];
    end
    if (rst) begin
      \$23  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$48 ) begin end
    \$24  = write_ptr_0;
    if (\$2 ) begin
      \$24  = \$3 [5:0];
    end
    if (rst) begin
      \$24  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$48 ) begin end
    \$25  = write_ptr_1;
    if (\$4 ) begin
      \$25  = \$5 [5:0];
    end
    if (rst) begin
      \$25  = 6'h00;
    end
  end
  assign input__0__payload = output__0__payload;
  assign input__1__payload = output__1__payload;
  assign \credit_in__payload[0]  = credit_in__payload[5:0];
  assign \credit_in__payload[1]  = credit_in__payload[11:6];
  assign \$1  = credit_in__valid;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_0_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$49  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_0_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$49 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_0_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$50  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$50 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$50 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_1_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$51  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_1_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$51 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_south_vc_1_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$52  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$52 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$52 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:832" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west (credit_in__valid, clk, rst, \port$216$0 , \port$234$0 , output__0__ready, output__1__ready, output__0__valid, input__0__ready, output__1__valid, input__1__ready, input__0__valid, input__1__valid, credit_in__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$53  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  reg [5:0] \$22 ;
  reg [5:0] \$23 ;
  reg [5:0] \$24 ;
  reg [5:0] \$25 ;
  wire [6:0] \$3 ;
  wire \$4 ;
  wire [6:0] \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  input [11:0] credit_in__payload;
  wire [11:0] credit_in__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:822" *)
  wire [5:0] \credit_in__payload[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit_in__valid;
  wire credit_in__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  wire input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  wire input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  wire [3:0] output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  input [2:0] \port$216$0 ;
  wire [2:0] \port$216$0 ;
  input [2:0] \port$234$0 ;
  wire [2:0] \port$234$0 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  reg [5:0] read_ptr_1 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_0 = 6'h00;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  reg [5:0] write_ptr_1 = 6'h00;
  assign \$2  = output__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__0__ready;
  assign \$3  = write_ptr_0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$4  = output__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:855" *) output__1__ready;
  assign \$5  = write_ptr_1 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *) 1'h1;
  assign \$6  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$7  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$8  = \$6  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$7 ;
  assign \$9  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$8 ;
  assign output__0__valid = input__0__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$9 ;
  assign \$10  = read_ptr_0[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[5];
  assign \$11  = read_ptr_0[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_0[4:0];
  assign \$12  = \$10  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$11 ;
  assign \$13  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$12 ;
  assign input__0__ready = output__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$13 ;
  assign \$14  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$15  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$16  = \$14  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$15 ;
  assign \$17  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$16 ;
  assign output__1__valid = input__1__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:851" *) \$17 ;
  assign \$18  = read_ptr_1[5] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[5];
  assign \$19  = read_ptr_1[4:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) write_ptr_1[4:0];
  assign \$20  = \$18  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:847" *) \$19 ;
  assign \$21  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$20 ;
  assign input__1__ready = output__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:852" *) \$21 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_0 <= \$22 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:834" *)
  always @(posedge clk)
    read_ptr_1 <= \$23 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_0 <= \$24 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:835" *)
  always @(posedge clk)
    write_ptr_1 <= \$25 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$53 ) begin end
    \$22  = read_ptr_0;
    if (\$1 ) begin
      \$22  = credit_in__payload[5:0];
    end
    if (rst) begin
      \$22  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$53 ) begin end
    \$23  = read_ptr_1;
    if (\$1 ) begin
      \$23  = credit_in__payload[11:6];
    end
    if (rst) begin
      \$23  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$53 ) begin end
    \$24  = write_ptr_0;
    if (\$2 ) begin
      \$24  = \$3 [5:0];
    end
    if (rst) begin
      \$24  = 6'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$53 ) begin end
    \$25  = write_ptr_1;
    if (\$4 ) begin
      \$25  = \$5 [5:0];
    end
    if (rst) begin
      \$25  = 6'h00;
    end
  end
  assign output__0__payload = { 1'h0, \port$216$0  };
  assign input__0__payload = { 1'h0, \port$216$0  };
  assign output__1__payload = { 1'h0, \port$234$0  };
  assign input__1__payload = { 1'h0, \port$234$0  };
  assign \credit_in__payload[0]  = credit_in__payload[5:0];
  assign \credit_in__payload[1]  = credit_in__payload[11:6];
  assign \$1  = credit_in__valid;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_0_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$54  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_0_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$54 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_0_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$55  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$55 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$55 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:999" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_1_arb (rst, input__0__valid, input__1__valid, input__2__valid, input__3__valid, input__4__valid, input__5__valid, input__6__valid, input__7__valid, output__ready, input__0__payload, input__1__payload, input__2__payload, input__3__payload, input__4__payload, input__5__payload, input__6__payload, input__7__payload, output__valid, output__payload, input__0__ready
, input__1__ready, input__2__ready, input__3__ready, input__4__ready, input__5__ready, input__6__ready, input__7__ready, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$56  = 0;
  reg \$1 ;
  wire \$10 ;
  reg \$11 ;
  reg \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* enum_base_type = "fsmState" *)
  (* enum_value_0 = "IDLE/0" *)
  (* enum_value_1 = "TRANSFER/1" *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  reg fsm_state = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  wire [2:0] grant_store;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1009" *)
  reg [2:0] granted;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  reg input__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  reg input__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__2__payload;
  wire input__2__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__2__ready;
  reg input__2__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__2__valid;
  wire input__2__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__3__payload;
  wire input__3__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__3__ready;
  reg input__3__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__3__valid;
  wire input__3__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__4__payload;
  wire input__4__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__4__ready;
  reg input__4__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__4__valid;
  wire input__4__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__5__payload;
  wire input__5__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__5__ready;
  reg input__5__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__5__valid;
  wire input__5__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__6__payload;
  wire input__6__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__6__ready;
  reg input__6__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__6__valid;
  wire input__6__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__7__payload;
  wire input__7__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__7__ready;
  reg input__7__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__7__valid;
  wire input__7__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  reg next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  output [3:0] output__payload;
  reg [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire \output__payload.last ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:992" *)
  wire [2:0] \output__payload.src ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  reg output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1010" *)
  reg transfer;
  assign \$3  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:485" *) fsm_state;
  assign \$6  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1023" *) requests;
  assign \$7  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__ready;
  assign \$8  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1029" *) output__payload[0];
  assign \$9  = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__ready;
  assign \$10  = \$9  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1038" *) output__payload[0];
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1039" *)
  always @(posedge clk)
    fsm_state <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:1004" *)
  \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_1_arb.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .grant_store(grant_store),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$1  = input__0__valid;
      3'h1:
          \$1  = input__1__valid;
      3'h2:
          \$1  = input__2__valid;
      3'h3:
          \$1  = input__3__valid;
      3'h4:
          \$1  = input__4__valid;
      3'h5:
          \$1  = input__5__valid;
      3'h6:
          \$1  = input__6__valid;
      3'h7:
          \$1  = input__7__valid;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    (* full_case = 32'd1 *)
    casez (granted)
      3'h0:
          \$2  = input__0__payload;
      3'h1:
          \$2  = input__1__payload;
      3'h2:
          \$2  = input__2__payload;
      3'h3:
          \$2  = input__3__payload;
      3'h4:
          \$2  = input__4__payload;
      3'h5:
          \$2  = input__5__payload;
      3'h6:
          \$2  = input__6__payload;
      3'h7:
          \$2  = input__7__payload;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    output__valid = 1'h0;
    if (transfer) begin
      output__valid = \$1 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    output__payload = 4'h0;
    if (transfer) begin
      output__payload[0] = \$2 ;
      output__payload[3:1] = granted;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__0__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            input__0__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__1__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            input__1__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__2__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            input__2__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__3__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            input__3__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__4__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            input__4__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__5__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            input__5__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__6__ready = 1'h0;
    if (transfer) begin
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            input__6__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    input__7__ready = 1'h0;
    if (transfer) begin
      (* full_case = 32'd1 *)
      casez (granted)
        3'h0:
            /* empty */;
        3'h1:
            /* empty */;
        3'h2:
            /* empty */;
        3'h3:
            /* empty */;
        3'h4:
            /* empty */;
        3'h5:
            /* empty */;
        3'h6:
            /* empty */;
        3'h7:
            input__7__ready = output__ready;
      endcase
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    next = 1'h0;
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            next = 1'h1;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    granted = 3'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            granted = grant;
          end
      1'h1:
          granted = grant_store;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    transfer = 1'h0;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$3 ) begin
            transfer = 1'h1;
          end
      1'h1:
          transfer = 1'h1;
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$56 ) begin end
    \$11  = fsm_state;
    (* full_case = 32'd1 *)
    casez (fsm_state)
      1'h0:
          if (\$6 ) begin
            (* full_case = 32'd1 *)
            if (\$8 ) begin
              \$11  = 1'h0;
            end else begin
              \$11  = 1'h1;
            end
          end
      1'h1:
          if (\$10 ) begin
            \$11  = 1'h0;
          end
    endcase
    if (rst) begin
      \$11  = 1'h0;
    end
  end
  assign \output__payload.last  = output__payload[0];
  assign \output__payload.src  = output__payload[3:1];
  assign requests[7] = input__7__valid;
  assign requests[6] = input__6__valid;
  assign requests[5] = input__5__valid;
  assign requests[4] = input__4__valid;
  assign requests[3] = input__3__valid;
  assign requests[2] = input__2__valid;
  assign requests[1] = input__1__valid;
  assign requests[0] = input__0__valid;
  assign \$5  = fsm_state;
endmodule

(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.RouterCrossbar.vc_allocator.credit_counter_tx_west_vc_1_arb.arbiter (rst, requests, next, grant, grant_store, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$57  = 0;
  reg [2:0] \$1 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output [2:0] grant;
  reg [2:0] grant;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  output [2:0] grant_store;
  reg [2:0] grant_store = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [7:0] requests;
  wire [7:0] requests;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$57 ) begin end
    grant = 3'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      3'h0:
        begin
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
        end
      3'h1:
        begin
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
        end
      3'h2:
        begin
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
        end
      3'h3:
        begin
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
        end
      3'h4:
        begin
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
        end
      3'h5:
        begin
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
        end
      3'h6:
        begin
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
          if (requests[7]) begin
            grant = 3'h7;
          end
        end
      3'h7:
        begin
          if (requests[7]) begin
            grant = 3'h7;
          end
          if (requests[6]) begin
            grant = 3'h6;
          end
          if (requests[5]) begin
            grant = 3'h5;
          end
          if (requests[4]) begin
            grant = 3'h4;
          end
          if (requests[3]) begin
            grant = 3'h3;
          end
          if (requests[2]) begin
            grant = 3'h2;
          end
          if (requests[1]) begin
            grant = 3'h1;
          end
          if (requests[0]) begin
            grant = 3'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$57 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 3'h0;
    end
  end
endmodule


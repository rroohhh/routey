

package multi_queue_credit_counter_tx_pkg;

endpackage

interface multi_queue_credit_counter_tx_in_stream_if import multi_queue_credit_counter_tx_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface multi_queue_credit_counter_tx_out_stream_if import multi_queue_credit_counter_tx_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface multi_queue_credit_counter_tx_credit_in_stream_if import multi_queue_credit_counter_tx_pkg::*;;
    logic [3: 0] payload[2];
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module multi_queue_credit_counter_tx import multi_queue_credit_counter_tx_pkg::*;
 (
    input wire clk,
    input wire rst,
    multi_queue_credit_counter_tx_in_stream_if.slave in[2],
    multi_queue_credit_counter_tx_out_stream_if.master out[2],
    multi_queue_credit_counter_tx_credit_in_stream_if.slave credit_in
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueCreditCounterTX
    \arq.MultiQueueCreditCounterTX  multi_queue_credit_counter_tx_internal (
        .clk,
        .rst,
        .input__0__payload(in[0].p),
        .input__0__valid(in[0].valid),
        .input__0__ready(in[0].ready),
        .input__1__payload(in[1].p),
        .input__1__valid(in[1].valid),
        .input__1__ready(in[1].ready),
        .output__0__payload(out[0].p),
        .output__0__valid(out[0].valid),
        .output__0__ready(out[0].ready),
        .output__1__payload(out[1].p),
        .output__1__valid(out[1].valid),
        .output__1__ready(out[1].ready),
        .credit_in__payload({<<4{credit_in.p}}),
        .credit_in__valid(credit_in.valid)
    );

    assign credit_in.ready = 1'd1;
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:741" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueCreditCounterTX (input__0__valid, input__1__payload, input__1__valid, output__0__ready, output__1__ready, credit_in__payload, credit_in__valid, clk, rst, input__0__ready, input__1__ready, output__0__payload, output__0__valid, output__1__payload, output__1__valid, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  reg [3:0] \$22 ;
  reg [3:0] \$23 ;
  reg [3:0] \$24 ;
  reg [3:0] \$25 ;
  wire [4:0] \$3 ;
  wire \$4 ;
  wire [4:0] \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:731" *)
  input [7:0] credit_in__payload;
  wire [7:0] credit_in__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:731" *)
  wire [3:0] \credit_in__payload[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:731" *)
  wire [3:0] \credit_in__payload[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input credit_in__valid;
  wire credit_in__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  wire input__0__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  wire input__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__0__payload;
  wire output__0__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__1__payload;
  wire output__1__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:743" *)
  reg [3:0] read_ptr_0 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:743" *)
  reg [3:0] read_ptr_1 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:744" *)
  reg [3:0] write_ptr_0 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:744" *)
  reg [3:0] write_ptr_1 = 4'h0;
  assign \$2  = output__0__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:764" *) output__0__ready;
  assign \$3  = write_ptr_0 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:765" *) 1'h1;
  assign \$4  = output__1__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:764" *) output__1__ready;
  assign \$5  = write_ptr_1 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:765" *) 1'h1;
  assign \$6  = read_ptr_0[3] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_0[3];
  assign \$7  = read_ptr_0[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_0[2:0];
  assign \$8  = \$6  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) \$7 ;
  assign \$9  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:760" *) \$8 ;
  assign output__0__valid = input__0__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:760" *) \$9 ;
  assign \$10  = read_ptr_0[3] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_0[3];
  assign \$11  = read_ptr_0[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_0[2:0];
  assign \$12  = \$10  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) \$11 ;
  assign \$13  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:761" *) \$12 ;
  assign input__0__ready = output__0__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:761" *) \$13 ;
  assign \$14  = read_ptr_1[3] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_1[3];
  assign \$15  = read_ptr_1[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_1[2:0];
  assign \$16  = \$14  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) \$15 ;
  assign \$17  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:760" *) \$16 ;
  assign output__1__valid = input__1__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:760" *) \$17 ;
  assign \$18  = read_ptr_1[3] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_1[3];
  assign \$19  = read_ptr_1[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) write_ptr_1[2:0];
  assign \$20  = \$18  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:756" *) \$19 ;
  assign \$21  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:761" *) \$20 ;
  assign input__1__ready = output__1__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:761" *) \$21 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:743" *)
  always @(posedge clk)
    read_ptr_0 <= \$22 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:743" *)
  always @(posedge clk)
    read_ptr_1 <= \$23 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:744" *)
  always @(posedge clk)
    write_ptr_0 <= \$24 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:744" *)
  always @(posedge clk)
    write_ptr_1 <= \$25 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$22  = read_ptr_0;
    if (\$1 ) begin
      \$22  = credit_in__payload[3:0];
    end
    if (rst) begin
      \$22  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$23  = read_ptr_1;
    if (\$1 ) begin
      \$23  = credit_in__payload[7:4];
    end
    if (rst) begin
      \$23  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$24  = write_ptr_0;
    if (\$2 ) begin
      \$24  = \$3 [3:0];
    end
    if (rst) begin
      \$24  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$25  = write_ptr_1;
    if (\$4 ) begin
      \$25  = \$5 [3:0];
    end
    if (rst) begin
      \$25  = 4'h0;
    end
  end
  assign output__0__payload = input__0__payload;
  assign output__1__payload = input__1__payload;
  assign \credit_in__payload[0]  = credit_in__payload[3:0];
  assign \credit_in__payload[1]  = credit_in__payload[7:4];
  assign \$1  = credit_in__valid;
endmodule




package arq_receiver_pkg;
typedef struct packed {
    logic p;
    logic [3: 0] seq;
} arq_payload;

typedef struct packed {
    logic seq_is_valid;
    logic is_nack;
    logic [3: 0] seq;
} ack;
endpackage

interface arq_receiver_out_stream_if import arq_receiver_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_payload_stream_if import arq_receiver_pkg::*;;
    arq_payload payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_receiver_ack_if import arq_receiver_pkg::*;;
    ack p;
    logic trigger;
    logic did_trigger;

    modport master (
        output p,
        output trigger,
        input did_trigger
    );
    modport slave (
        input p,
        input trigger,
        output did_trigger
    );
    modport monitor (
        input p,
        input trigger,
        input did_trigger
    );
endinterface

module arq_receiver import arq_receiver_pkg::*;
 (
    input wire clk,
    input wire rst,
    input wire logic input_error,
    arq_receiver_out_stream_if.master out,
    arq_payload_stream_if.slave in,
    arq_receiver_ack_if.master ack
);
    // connect_rpc -exec amaranth-rpc yosys arq.ArqReceiver
    \arq.ArqReceiver  arq_receiver_internal (
        .clk,
        .rst,
        .input_error(input_error),
        .output__payload(out.p),
        .output__valid(out.valid),
        .output__ready(out.ready),
        .input__payload(in.p),
        .input__valid(in.valid),
        .input__ready(in.ready),
        .ack__p(ack.p),
        .ack__trigger(ack.trigger),
        .ack__did_trigger(ack.did_trigger)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:297" *)
(* generator = "Amaranth" *)
module \arq.ArqReceiver (output__ready, input__payload, input__valid, ack__did_trigger, clk, rst, output__payload, output__valid, input__ready, ack__p, ack__trigger, input_error);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire [4:0] \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire [5:0] \$20 ;
  wire \$21 ;
  wire \$22 ;
  wire \$23 ;
  wire \$24 ;
  wire \$25 ;
  wire [1:0] \$26 ;
  reg \$27 ;
  reg [3:0] \$28 ;
  reg [4:0] \$29 ;
  wire \$3 ;
  reg \$30 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:46" *)
  input ack__did_trigger;
  wire ack__did_trigger;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:289" *)
  output [5:0] ack__p;
  reg [5:0] ack__p;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:289" *)
  wire \ack__p.is_nack ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:289" *)
  wire [3:0] \ack__p.seq ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:289" *)
  wire \ack__p.seq_is_valid ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:45" *)
  output ack__trigger;
  reg ack__trigger;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:301" *)
  wire [3:0] expected_seq;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:289" *)
  input [4:0] input__payload;
  wire [4:0] input__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:289" *)
  wire \input__payload.p ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:289" *)
  wire [3:0] \input__payload.seq ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:290" *)
  input input_error;
  wire input_error;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:299" *)
  reg [3:0] last_seq = 4'hf;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:300" *)
  reg last_seq_valid = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__payload;
  wire output__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:336" *)
  reg [4:0] timeout_counter = 5'h00;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:329" *)
  reg word_counter = 1'h0;
  assign \$1  = last_seq + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:302" *) 1'h1;
  assign \$2  = input__payload[3:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$1 [3:0];
  assign \$3  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$2 ;
  assign \$4  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:311" *) \$3 ;
  assign \$5  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:311" *) \$4 ;
  assign input__ready = output__ready | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:311" *) \$5 ;
  assign \$6  = input__payload[3:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$1 [3:0];
  assign output__valid = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$6 ;
  assign \$7  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:338" *) word_counter;
  assign \$8  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:341" *) timeout_counter;
  assign \$9  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:303" *) input__ready;
  assign \$10  = input__payload[3:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$1 [3:0];
  assign \$11  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$10 ;
  assign \$12  = \$9  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:348" *) \$11 ;
  assign \$14  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:303" *) input__ready;
  assign \$15  = input__payload[3:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$1 [3:0];
  assign \$16  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$15 ;
  assign \$17  = \$14  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:306" *) \$16 ;
  assign \$18  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:338" *) word_counter;
  assign \$19  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:341" *) timeout_counter;
  assign \$20  = timeout_counter - (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:342" *) 1'h1;
  assign \$21  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:303" *) input__ready;
  assign \$22  = input__payload[3:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$1 [3:0];
  assign \$23  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:305" *) \$22 ;
  assign \$24  = \$21  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:348" *) \$23 ;
  assign \$26  = word_counter + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:353" *) 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:300" *)
  always @(posedge clk)
    last_seq_valid <= \$27 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:299" *)
  always @(posedge clk)
    last_seq <= \$28 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:336" *)
  always @(posedge clk)
    timeout_counter <= \$29 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:329" *)
  always @(posedge clk)
    word_counter <= \$30 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    ack__p[4] = 1'h0;
    (* full_case = 32'd1 *)
    if (\$7 ) begin
    end else begin
      (* full_case = 32'd1 *)
      if (\$8 ) begin
      end else begin
        ack__p[4] = 1'h0;
      end
    end
    if (\$12 ) begin
      if (\$13 ) begin
        ack__p[4] = 1'h0;
      end
    end
    if (input_error) begin
      ack__p[4] = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    ack__trigger = 1'h0;
    (* full_case = 32'd1 *)
    if (\$7 ) begin
    end else begin
      (* full_case = 32'd1 *)
      if (\$8 ) begin
      end else begin
        ack__trigger = 1'h1;
      end
    end
    if (\$12 ) begin
      if (\$13 ) begin
        ack__trigger = 1'h1;
      end
    end
    if (input_error) begin
      ack__trigger = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$27  = last_seq_valid;
    if (\$17 ) begin
      \$27  = 1'h1;
    end
    if (rst) begin
      \$27  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$28  = last_seq;
    if (\$17 ) begin
      \$28  = input__payload[3:0];
    end
    if (rst) begin
      \$28  = 4'hf;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (\$18 ) begin
      \$29  = 5'h10;
    end else begin
      (* full_case = 32'd1 *)
      if (\$19 ) begin
        \$29  = \$20 [4:0];
      end else begin
        \$29  = 5'h10;
      end
    end
    if (rst) begin
      \$29  = 5'h00;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$30  = word_counter;
    if (\$24 ) begin
      (* full_case = 32'd1 *)
      if (\$25 ) begin
        \$30  = 1'h0;
      end else begin
        \$30  = \$26 [0];
      end
    end
    if (ack__did_trigger) begin
      \$30  = 1'h0;
    end
    if (rst) begin
      \$30  = 1'h0;
    end
  end
  assign expected_seq = \$1 [3:0];
  assign output__payload = input__payload[4];
  assign \input__payload.seq  = input__payload[3:0];
  assign \input__payload.p  = input__payload[4];
  assign \ack__p.seq  = ack__p[3:0];
  assign \ack__p.is_nack  = ack__p[4];
  assign \ack__p.seq_is_valid  = ack__p[5];
  always @*
    ack__p[5] = last_seq_valid;
  always @*
    ack__p[3:0] = last_seq;
  assign \$13  = word_counter;
  assign \$25  = word_counter;
endmodule




package multi_queue_fifo_reader_pkg;

endpackage

interface multi_queue_fifo_reader_in_stream_if import multi_queue_fifo_reader_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface multi_queue_fifo_reader_out_stream_if import multi_queue_fifo_reader_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module multi_queue_fifo_reader import multi_queue_fifo_reader_pkg::*;
 (
    input wire clk,
    input wire rst,
    multi_queue_fifo_reader_in_stream_if.slave in[2],
    multi_queue_fifo_reader_out_stream_if.master out[2]
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueFifoReader
    \arq.MultiQueueFifoReader  multi_queue_fifo_reader_internal (
        .clk,
        .rst,
        .input__0__payload(in[0].p),
        .input__0__valid(in[0].valid),
        .input__0__ready(in[0].ready),
        .input__1__payload(in[1].p),
        .input__1__valid(in[1].valid),
        .input__1__ready(in[1].ready),
        .output__0__payload(out[0].p),
        .output__0__valid(out[0].valid),
        .output__0__ready(out[0].ready),
        .output__1__payload(out[1].p),
        .output__1__valid(out[1].valid),
        .output__1__ready(out[1].ready)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:936" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueFifoReader (input__0__valid, input__1__payload, input__1__valid, output__0__ready, output__1__ready, clk, rst, input__0__ready, input__1__ready, output__0__payload, output__0__valid, output__1__payload, output__1__valid, input__0__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  reg \$19 ;
  wire \$2 ;
  reg \$20 ;
  wire \$3 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  wire grant;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__0__payload;
  wire input__0__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__0__ready;
  wire input__0__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__0__valid;
  wire input__0__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  input input__1__payload;
  wire input__1__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__1__ready;
  wire input__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__1__valid;
  wire input__1__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  wire next;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__0__payload;
  wire output__0__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__1__payload;
  wire output__1__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:944" *)
  reg ready_outstanding_0 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:944" *)
  reg ready_outstanding_1 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  wire [1:0] requests;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  assign next = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:939" *) requests;
  assign \$1  = input__0__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:950" *) output__0__ready;
  assign \$2  = \$1  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:950" *) ready_outstanding_0;
  assign \$3  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:951" *) requests;
  assign \$4  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:951" *) grant;
  assign input__0__ready = \$3  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:951" *) \$4 ;
  assign \$5  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:952" *) ready_outstanding_0;
  assign output__0__valid = input__0__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:952" *) \$5 ;
  assign \$6  = input__1__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:950" *) output__1__ready;
  assign \$7  = \$6  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:950" *) ready_outstanding_1;
  assign \$8  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:951" *) requests;
  assign input__1__ready = \$8  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:951" *) \$9 ;
  assign \$10  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:952" *) ready_outstanding_1;
  assign output__1__valid = input__1__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:952" *) \$10 ;
  assign \$11  = output__0__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:956" *) output__0__ready;
  assign \$12  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:956" *) input__0__ready;
  assign \$13  = \$11  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:956" *) \$12 ;
  assign \$14  = ready_outstanding_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:959" *) input__0__ready;
  assign \$15  = output__1__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:956" *) output__1__ready;
  assign \$16  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:956" *) input__1__ready;
  assign \$17  = \$15  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:956" *) \$16 ;
  assign \$18  = ready_outstanding_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:959" *) input__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:944" *)
  always @(posedge clk)
    ready_outstanding_0 <= \$19 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:944" *)
  always @(posedge clk)
    ready_outstanding_1 <= \$20 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:938" *)
  \arq.MultiQueueFifoReader.arbiter  arbiter (
    .clk(clk),
    .grant(grant),
    .next(next),
    .requests(requests),
    .rst(rst)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$19  = ready_outstanding_0;
    if (\$13 ) begin
      \$19  = 1'h1;
    end
    if (\$14 ) begin
      \$19  = 1'h0;
    end
    if (rst) begin
      \$19  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$20  = ready_outstanding_1;
    if (\$17 ) begin
      \$20  = 1'h1;
    end
    if (\$18 ) begin
      \$20  = 1'h0;
    end
    if (rst) begin
      \$20  = 1'h0;
    end
  end
  assign output__0__payload = input__0__payload;
  assign output__1__payload = input__1__payload;
  assign requests[1] = \$7 ;
  assign requests[0] = \$2 ;
  assign \$9  = grant;
endmodule

(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:19" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueFifoReader.arbiter (rst, next, requests, grant, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$2  = 0;
  reg \$1 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:15" *)
  output grant;
  reg grant;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  reg grant_store = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:13" *)
  input next;
  wire next;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:12" *)
  input [1:0] requests;
  wire [1:0] requests;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/round_robin_arbiter.py:14" *)
  always @(posedge clk)
    grant_store <= \$1 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    grant = 1'h0;
    (* full_case = 32'd1 *)
    casez (grant_store)
      1'h0:
        begin
          if (requests[0]) begin
            grant = 1'h0;
          end
          if (requests[1]) begin
            grant = 1'h1;
          end
        end
      1'h1:
        begin
          if (requests[1]) begin
            grant = 1'h1;
          end
          if (requests[0]) begin
            grant = 1'h0;
          end
        end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    \$1  = grant_store;
    if (next) begin
      \$1  = grant;
    end
    if (rst) begin
      \$1  = 1'h0;
    end
  end
endmodule


package flit_tag;
typedef enum logic [2: 0] {
    START = 0,
    TAIL = 1,
    PAYLOAD = 2,
    START_AND_END = 3,
    ARQ_ACK = 4
} flit_tag;
endpackage

package cardinal_port;
typedef enum logic [2: 0] {
    LOCAL = 0,
    NORTH = 1,
    SOUTH = 2,
    EAST = 3,
    WEST = 4
} cardinal_port;
endpackage

package input_channel_pkg;
import flit_tag::flit_tag;
import cardinal_port::cardinal_port;
export flit_tag::flit_tag;
export cardinal_port::cardinal_port;
typedef logic [5: 0][1:0] flit_arqack_credit;

typedef struct packed {
    logic [59: 0] payload;
    logic is_nack;
    logic seq_is_valid;
    flit_arqack_credit credit;
} flit_arqack;

typedef struct packed {
    logic [6: 0] y;
    logic [6: 0] x;
} coordinate;

typedef struct packed {
    coordinate target;
} routing_target;

typedef struct packed {
    logic [59: 0] payload;
    routing_target target;
} flit_start_and_end;

typedef struct packed {
    logic [73: 0] payload;
} flit_payload;

typedef struct packed {
    logic [73: 0] payload;
} flit_tail;

typedef struct packed {
    logic [59: 0] payload;
    routing_target target;
} flit_start;

typedef union packed {
    flit_arqack arq_ack;
    flit_start_and_end start_and_end;
    flit_payload payload;
    flit_tail tail;
    flit_start start;
} flit_data;

typedef struct packed {
    flit_data data;
    flit_tag tag;
} flit;

typedef struct packed {
    logic vc_id;
    cardinal_port port;
} port;

typedef struct packed {
    port target;
    logic last;
    flit flit;
} routed_flit;
endpackage

interface flit_stream_if import input_channel_pkg::*;;
    flit payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface routed_flit_stream_if import input_channel_pkg::*;;
    routed_flit payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface input_channel_cfg_if import input_channel_pkg::*;;
    logic [31: 0] invalid_flit_ctr;

    modport master (
        input invalid_flit_ctr
    );
    modport slave (
        output invalid_flit_ctr
    );
    modport monitor (
        input invalid_flit_ctr
    );
endinterface

interface input_channel_route_computer_cfg_if import input_channel_pkg::*;;
    coordinate position;

    modport master (
        output position
    );
    modport slave (
        input position
    );
    modport monitor (
        input position
    );
endinterface

module input_channel import input_channel_pkg::*;
 (
    input wire clk,
    input wire rst,
    flit_stream_if.slave flit_in,
    routed_flit_stream_if.master flit_out,
    input_channel_cfg_if.slave cfg,
    input_channel_route_computer_cfg_if.slave route_computer_cfg
);
    // connect_rpc -exec amaranth-rpc yosys memory_mapped_router.InputChannel
    \memory_mapped_router.InputChannel  input_channel_internal (
        .clk,
        .rst,
        .flit_in__payload(flit_in.p),
        .flit_in__valid(flit_in.valid),
        .flit_in__ready(flit_in.ready),
        .flit_out__payload(flit_out.p),
        .flit_out__valid(flit_out.valid),
        .flit_out__ready(flit_out.ready),
        .cfg__invalid_flit_ctr(cfg.invalid_flit_ctr),
        .route_computer_cfg__position(route_computer_cfg.position)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:223" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.InputChannel (flit_in__valid, flit_out__ready, route_computer_cfg__position, clk, rst, flit_in__ready, flit_out__payload, flit_out__valid, cfg__invalid_flit_ctr, flit_in__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  wire \$22 ;
  wire \$23 ;
  wire \$24 ;
  wire \$25 ;
  reg \$26 ;
  reg \$27 ;
  reg \$28 ;
  wire \$3 ;
  wire [13:0] \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:205" *)
  output [31:0] cfg__invalid_flit_ctr;
  wire [31:0] cfg__invalid_flit_ctr;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] cfg__position;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \cfg__position.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \cfg__position.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  input [76:0] flit_in__payload;
  wire [76:0] flit_in__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output flit_in__ready;
  wire flit_in__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input flit_in__valid;
  wire flit_in__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:217" *)
  output [81:0] flit_out__payload;
  wire [81:0] flit_out__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:217" *)
  wire \flit_out__payload.last ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:217" *)
  wire [3:0] \flit_out__payload.target ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:217" *)
  wire [2:0] \flit_out__payload.target.port ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:217" *)
  wire \flit_out__payload.target.vc_id ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input flit_out__ready;
  wire flit_out__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output flit_out__valid;
  wire flit_out__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [14:0] input__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \input__payload.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \input__payload.target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \input__payload.target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \input__payload.target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire \input__payload.vc ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire input__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  reg input__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:233" *)
  reg next_flit_in_has_routing = 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:277" *)
  reg next_flit_out_has_routing = 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [76:0] r_stream__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [17:0] \r_stream__payload$29 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \r_stream__payload$29.new_target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \r_stream__payload$29.new_target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \r_stream__payload$29.new_target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \r_stream__payload$29.new_target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [3:0] \r_stream__payload$29.port ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [2:0] \r_stream__payload$29.port.port ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire \r_stream__payload$29.port.vc_id ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire r_stream__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \r_stream__ready$32 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire r_stream__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \r_stream__valid$31 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [17:0] result__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \result__payload.new_target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \result__payload.new_target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \result__payload.new_target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \result__payload.new_target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [3:0] \result__payload.port ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [2:0] \result__payload.port.port ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire \result__payload.port.vc_id ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire result__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire result__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  input [13:0] route_computer_cfg__position;
  wire [13:0] route_computer_cfg__position;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:217" *)
  wire [6:0] \route_computer_cfg__position.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:217" *)
  wire [6:0] \route_computer_cfg__position.y ;
  (* enum_base_type = "route_computer_fsmState" *)
  (* enum_value_0 = "idle/0" *)
  (* enum_value_1 = "wait_for_new/1" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:265" *)
  reg route_computer_fsm_state = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:237" *)
  reg route_computer_stall;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [76:0] w_stream__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [17:0] \w_stream__payload$20 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \w_stream__payload$20.new_target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \w_stream__payload$20.new_target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \w_stream__payload$20.new_target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \w_stream__payload$20.new_target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [3:0] \w_stream__payload$20.port ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [2:0] \w_stream__payload$20.port.port ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire \w_stream__payload$20.port.vc_id ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire w_stream__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire \w_stream__ready$23 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire w_stream__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire \w_stream__valid$24 ;
  assign \$1  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:241" *) route_computer_stall;
  assign flit_in__ready = w_stream__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:241" *) \$1 ;
  assign \$2  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:242" *) route_computer_stall;
  assign w_stream__valid = flit_in__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:242" *) \$2 ;
  assign \$3  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:257" *) input__ready;
  assign r_stream__ready = flit_out__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:283" *) flit_out__valid;
  assign \$4  = next_flit_out_has_routing ? (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:285" *) \r_stream__payload$29 [13:0] : r_stream__payload[16:3];
  assign \$5  = r_stream__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$6  = r_stream__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$7  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$6 , \$5  };
  assign flit_out__valid = r_stream__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:290" *) \r_stream__valid$31 ;
  assign \$8  = flit_out__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:291" *) flit_out__valid;
  assign \$9  = flit_out__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$10  = flit_out__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$11  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$10 , \$9  };
  assign \r_stream__ready$32  = \$8  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:291" *) \$11 ;
  assign \$12  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_dsl.py:486" *) route_computer_fsm_state;
  assign \$14  = flit_in__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:234" *) flit_in__ready;
  assign \$15  = flit_in__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$16  = flit_in__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$17  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$16 , \$15  };
  assign \$18  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:261" *) input__ready;
  assign \$19  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:261" *) w_stream__ready;
  assign \$20  = \$18  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:261" *) \$19 ;
  assign \$21  = w_stream__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:264" *) w_stream__ready;
  assign \$22  = flit_out__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:278" *) flit_out__ready;
  assign \$23  = flit_out__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 2'h3;
  assign \$24  = flit_out__payload[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1315" *) 1'h1;
  assign \$25  = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ast.py:1321" *) { \$24 , \$23  };
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:233" *)
  always @(posedge clk)
    next_flit_in_has_routing <= \$26 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:265" *)
  always @(posedge clk)
    route_computer_fsm_state <= \$27 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:277" *)
  always @(posedge clk)
    next_flit_out_has_routing <= \$28 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:229" *)
  \memory_mapped_router.InputChannel.input_fifo  input_fifo (
    .clk(clk),
    .r_en(r_stream__ready),
    .r_stream__payload(r_stream__payload),
    .r_stream__valid(r_stream__valid),
    .rst(rst),
    .w_data(flit_in__payload),
    .w_en(w_stream__valid),
    .w_stream__ready(w_stream__ready)
  );
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  \memory_mapped_router.InputChannel.route_computer  route_computer (
    .cfg__position(route_computer_cfg__position),
    .input__payload(input__payload),
    .input__ready(input__ready),
    .result__payload(\w_stream__payload$20 ),
    .result__valid(input__valid)
  );
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:267" *)
  \memory_mapped_router.InputChannel.route_result_fifo  route_result_fifo (
    .clk(clk),
    .r_en(\r_stream__ready$32 ),
    .r_stream__payload(\r_stream__payload$29 ),
    .r_stream__valid(\r_stream__valid$31 ),
    .rst(rst),
    .w_data(\w_stream__payload$20 ),
    .w_en(input__valid),
    .w_stream__ready(input__ready)
  );
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    input__valid = 1'h0;
    casez (route_computer_fsm_state)
      1'h0:
          if (next_flit_in_has_routing) begin
            input__valid = flit_in__valid;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    route_computer_stall = 1'h0;
    casez (route_computer_fsm_state)
      1'h0:
          if (next_flit_in_has_routing) begin
            route_computer_stall = \$3 ;
          end
    endcase
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$26  = next_flit_in_has_routing;
    if (\$14 ) begin
      \$26  = \$17 ;
    end
    if (rst) begin
      \$26  = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$27  = route_computer_fsm_state;
    (* full_case = 32'd1 *)
    casez (route_computer_fsm_state)
      1'h0:
          if (next_flit_in_has_routing) begin
            if (\$20 ) begin
              \$27  = 1'h1;
            end
          end
      1'h1:
          if (\$21 ) begin
            \$27  = 1'h0;
          end
    endcase
    if (rst) begin
      \$27  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$28  = next_flit_out_has_routing;
    if (\$22 ) begin
      \$28  = \$25 ;
    end
    if (rst) begin
      \$28  = 1'h1;
    end
  end
  assign cfg__position = route_computer_cfg__position;
  assign w_stream__payload = flit_in__payload;
  assign result__payload = \w_stream__payload$20 ;
  assign result__ready = input__ready;
  assign \w_stream__ready$23  = input__ready;
  assign \w_stream__valid$24  = input__valid;
  assign result__valid = input__valid;
  assign cfg__invalid_flit_ctr = 32'd0;
  assign \flit_out__payload.last  = flit_out__payload[77];
  assign \flit_out__payload.target  = flit_out__payload[81:78];
  assign \flit_out__payload.target.port  = flit_out__payload[80:78];
  assign \flit_out__payload.target.vc_id  = flit_out__payload[81];
  assign \route_computer_cfg__position.x  = route_computer_cfg__position[6:0];
  assign \route_computer_cfg__position.y  = route_computer_cfg__position[13:7];
  assign \cfg__position.x  = route_computer_cfg__position[6:0];
  assign \cfg__position.y  = route_computer_cfg__position[13:7];
  assign \input__payload.vc  = input__payload[0];
  assign \input__payload.target  = input__payload[14:1];
  assign \input__payload.target.target  = input__payload[14:1];
  assign \input__payload.target.target.x  = input__payload[7:1];
  assign \input__payload.target.target.y  = input__payload[14:8];
  assign \w_stream__payload$20.new_target  = \w_stream__payload$20 [13:0];
  assign \w_stream__payload$20.new_target.target  = \w_stream__payload$20 [13:0];
  assign \w_stream__payload$20.new_target.target.x  = \w_stream__payload$20 [6:0];
  assign \w_stream__payload$20.new_target.target.y  = \w_stream__payload$20 [13:7];
  assign \w_stream__payload$20.port  = \w_stream__payload$20 [17:14];
  assign \w_stream__payload$20.port.port  = \w_stream__payload$20 [16:14];
  assign \w_stream__payload$20.port.vc_id  = \w_stream__payload$20 [17];
  assign \result__payload.new_target  = \w_stream__payload$20 [13:0];
  assign \result__payload.new_target.target  = \w_stream__payload$20 [13:0];
  assign \result__payload.new_target.target.x  = \w_stream__payload$20 [6:0];
  assign \result__payload.new_target.target.y  = \w_stream__payload$20 [13:7];
  assign \result__payload.port  = \w_stream__payload$20 [17:14];
  assign \result__payload.port.port  = \w_stream__payload$20 [16:14];
  assign \result__payload.port.vc_id  = \w_stream__payload$20 [17];
  assign \r_stream__payload$29.new_target  = \r_stream__payload$29 [13:0];
  assign \r_stream__payload$29.new_target.target  = \r_stream__payload$29 [13:0];
  assign \r_stream__payload$29.new_target.target.x  = \r_stream__payload$29 [6:0];
  assign \r_stream__payload$29.new_target.target.y  = \r_stream__payload$29 [13:7];
  assign \r_stream__payload$29.port  = \r_stream__payload$29 [17:14];
  assign \r_stream__payload$29.port.port  = \r_stream__payload$29 [16:14];
  assign \r_stream__payload$29.port.vc_id  = \r_stream__payload$29 [17];
  assign flit_out__payload[77] = \$7 ;
  assign flit_out__payload[81:78] = \r_stream__payload$29 [17:14];
  assign flit_out__payload[2:0] = r_stream__payload[2:0];
  assign flit_out__payload[76:17] = r_stream__payload[76:17];
  assign flit_out__payload[16:3] = \$4 ;
  assign input__payload[0] = 1'h0;
  assign input__payload[14:1] = flit_in__payload[16:3];
  assign \$13  = route_computer_fsm_state;
endmodule

(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:36" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.InputChannel.input_fifo (clk, rst, w_en, r_en, w_stream__ready, r_stream__valid, r_stream__payload, w_data);
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:92" *)
  wire [76:0] r_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input r_en;
  wire r_en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:93" *)
  wire r_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:92" *)
  output [76:0] r_stream__payload;
  wire [76:0] r_stream__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire r_stream__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:93" *)
  output r_stream__valid;
  wire r_stream__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  input [76:0] w_data;
  wire [76:0] w_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input w_en;
  wire w_en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:88" *)
  wire w_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [76:0] w_stream__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:88" *)
  output w_stream__ready;
  wire w_stream__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire w_stream__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:40" *)
  \memory_mapped_router.InputChannel.input_fifo.fifo  fifo (
    .clk(clk),
    .r_data(r_stream__payload),
    .r_en(r_en),
    .r_rdy(r_stream__valid),
    .rst(rst),
    .w_en(w_en),
    .w_port__data(w_data),
    .w_rdy(w_stream__ready)
  );
  assign r_data = r_stream__payload;
  assign r_stream__ready = r_en;
  assign r_rdy = r_stream__valid;
  assign w_stream__payload = w_data;
  assign w_rdy = w_stream__ready;
  assign w_stream__valid = w_en;
endmodule

(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:144" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.InputChannel.input_fifo.fifo (clk, rst, w_en, r_en, w_rdy, r_rdy, r_data, w_port__data);
  reg \$auto$verilog_backend.cc:2355:dump_module$2  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire [2:0] \$14 ;
  reg \$15 ;
  reg \$16 ;
  reg [1:0] \$17 ;
  wire [1:0] \$2 ;
  wire \$3 ;
  wire [1:0] \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire [2:0] \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* init = 1'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:166" *)
  wire consume;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:141" *)
  reg [1:0] level = 2'h0;
  (* init = 1'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:165" *)
  wire produce;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:241" *)
  output [76:0] r_data;
  wire [76:0] r_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:94" *)
  input r_en;
  wire r_en;
  (* init = 2'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:95" *)
  wire [1:0] r_level;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:240" *)
  reg r_port__addr = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:241" *)
  wire [76:0] r_port__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:93" *)
  output r_rdy;
  wire r_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:87" *)
  wire [76:0] w_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:89" *)
  input w_en;
  wire w_en;
  (* init = 2'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:90" *)
  wire [1:0] w_level;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:401" *)
  reg w_port__addr = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:87" *)
  input [76:0] w_port__data;
  wire [76:0] w_port__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:400" *)
  wire w_port__en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:88" *)
  output w_rdy;
  wire w_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:162" *)
  reg [76:0] storage [1:0];
  initial begin
    storage[0] = 77'h00000000000000000000;
    storage[1] = 77'h00000000000000000000;
  end
  always @(posedge clk) begin
    if (w_port__en)
      storage[w_port__addr] <= w_port__data;
  end
  assign r_data = storage[r_port__addr];
  assign w_rdy = level != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:153" *) 2'h2;
  assign r_rdy = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:154" *) level;
  assign w_port__en = w_en & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:171" *) w_rdy;
  assign \$1  = w_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:160" *) w_en;
  assign \$2  = w_port__addr + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:116" *) 1'h1;
  assign \$3  = r_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:159" *) r_en;
  assign \$4  = r_port__addr + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:116" *) 1'h1;
  assign \$5  = w_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:160" *) w_en;
  assign \$6  = r_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:159" *) r_en;
  assign \$7  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:183" *) \$6 ;
  assign \$8  = \$5  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:183" *) \$7 ;
  assign \$9  = level + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:184" *) 1'h1;
  assign \$10  = r_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:159" *) r_en;
  assign \$11  = w_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:160" *) w_en;
  assign \$12  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:185" *) \$11 ;
  assign \$13  = \$10  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:185" *) \$12 ;
  assign \$14  = level - (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:186" *) 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:165" *)
  always @(posedge clk)
    w_port__addr <= \$15 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:166" *)
  always @(posedge clk)
    r_port__addr <= \$16 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:141" *)
  always @(posedge clk)
    level <= \$17 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    \$15  = w_port__addr;
    if (\$1 ) begin
      \$15  = \$2 [0];
    end
    if (rst) begin
      \$15  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    \$16  = r_port__addr;
    if (\$3 ) begin
      \$16  = \$4 [0];
    end
    if (rst) begin
      \$16  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$2 ) begin end
    \$17  = level;
    if (\$8 ) begin
      \$17  = \$9 [1:0];
    end
    if (\$13 ) begin
      \$17  = \$14 [1:0];
    end
    if (rst) begin
      \$17  = 2'h0;
    end
  end
  assign w_level = level;
  assign r_level = level;
  assign produce = w_port__addr;
  assign w_data = w_port__data;
  assign consume = r_port__addr;
  assign r_port__data = r_data;
endmodule

(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:170" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.InputChannel.route_computer (input__ready, input__payload, result__valid, result__payload, cfg__position);
  reg \$auto$verilog_backend.cc:2355:dump_module$3  = 0;
  wire \$1 ;
  wire \$2 ;
  wire \$3 ;
  wire [2:0] \$4 ;
  wire \$5 ;
  wire [2:0] \$6 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  input [13:0] cfg__position;
  wire [13:0] cfg__position;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \cfg__position.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \cfg__position.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  input [14:0] input__payload;
  wire [14:0] input__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \input__payload.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \input__payload.target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \input__payload.target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \input__payload.target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire \input__payload.vc ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input input__ready;
  wire input__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire input__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  output [17:0] result__payload;
  reg [17:0] result__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \result__payload.new_target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [13:0] \result__payload.new_target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \result__payload.new_target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [6:0] \result__payload.new_target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [3:0] \result__payload.port ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire [2:0] \result__payload.port.port ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:224" *)
  wire \result__payload.port.vc_id ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire result__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input result__valid;
  wire result__valid;
  assign \$4  = \$3  ? (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:186" *) 3'h3 : 3'h4;
  assign \$5  = input__payload[14:8] > (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:188" *) cfg__position[13:7];
  assign \$6  = \$5  ? (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:188" *) 3'h2 : 3'h1;
  assign \$1  = input__payload[7:1] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:185" *) cfg__position[6:0];
  assign \$2  = input__payload[14:8] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:187" *) cfg__position[13:7];
  assign \$3  = input__payload[7:1] > (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:186" *) cfg__position[6:0];
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$3 ) begin end
    (* full_case = 32'd1 *)
    if (\$1 ) begin
      result__payload[16:14] = \$4 ;
    end else if (\$2 ) begin
      result__payload[16:14] = \$6 ;
    end else begin
      result__payload[16:14] = 3'h0;
    end
  end
  assign result__ready = input__ready;
  assign input__valid = result__valid;
  assign \result__payload.new_target  = result__payload[13:0];
  assign \result__payload.new_target.target  = result__payload[13:0];
  assign \result__payload.new_target.target.x  = result__payload[6:0];
  assign \result__payload.new_target.target.y  = result__payload[13:7];
  assign \result__payload.port  = result__payload[17:14];
  assign \result__payload.port.port  = result__payload[16:14];
  assign \result__payload.port.vc_id  = result__payload[17];
  assign \input__payload.vc  = input__payload[0];
  assign \input__payload.target  = input__payload[14:1];
  assign \input__payload.target.target  = input__payload[14:1];
  assign \input__payload.target.target.x  = input__payload[7:1];
  assign \input__payload.target.target.y  = input__payload[14:8];
  assign \cfg__position.x  = cfg__position[6:0];
  assign \cfg__position.y  = cfg__position[13:7];
  always @*
    result__payload[17] = input__payload[0];
  always @*
    result__payload[13:0] = input__payload[14:1];
endmodule

(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:36" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.InputChannel.route_result_fifo (rst, r_en, w_stream__ready, r_stream__valid, r_stream__payload, w_en, w_data, clk);
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:92" *)
  wire [17:0] r_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input r_en;
  wire r_en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:93" *)
  wire r_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:92" *)
  output [17:0] r_stream__payload;
  wire [17:0] r_stream__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \r_stream__payload.new_target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \r_stream__payload.new_target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \r_stream__payload.new_target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \r_stream__payload.new_target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [3:0] \r_stream__payload.port ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [2:0] \r_stream__payload.port.port ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire \r_stream__payload.port.vc_id ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  wire r_stream__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:93" *)
  output r_stream__valid;
  wire r_stream__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  input [17:0] w_data;
  wire [17:0] w_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input w_en;
  wire w_en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:88" *)
  wire w_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [17:0] w_stream__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \w_stream__payload.new_target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [13:0] \w_stream__payload.new_target.target ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \w_stream__payload.new_target.target.x ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [6:0] \w_stream__payload.new_target.target.y ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [3:0] \w_stream__payload.port ;
  (* enum_base_type = "CardinalPort" *)
  (* enum_value_000 = "local" *)
  (* enum_value_001 = "north" *)
  (* enum_value_010 = "south" *)
  (* enum_value_011 = "east" *)
  (* enum_value_100 = "west" *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire [2:0] \w_stream__payload.port.port ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:29" *)
  wire \w_stream__payload.port.vc_id ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:88" *)
  output w_stream__ready;
  wire w_stream__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  wire w_stream__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/memory_mapped_router.py:40" *)
  \memory_mapped_router.InputChannel.route_result_fifo.fifo  fifo (
    .clk(clk),
    .r_data(r_stream__payload),
    .r_en(r_en),
    .r_rdy(r_stream__valid),
    .rst(rst),
    .w_en(w_en),
    .w_port__data(w_data),
    .w_rdy(w_stream__ready)
  );
  assign r_data = r_stream__payload;
  assign r_stream__ready = r_en;
  assign r_rdy = r_stream__valid;
  assign w_stream__payload = w_data;
  assign w_rdy = w_stream__ready;
  assign w_stream__valid = w_en;
  assign \r_stream__payload.new_target  = r_stream__payload[13:0];
  assign \r_stream__payload.new_target.target  = r_stream__payload[13:0];
  assign \r_stream__payload.new_target.target.x  = r_stream__payload[6:0];
  assign \r_stream__payload.new_target.target.y  = r_stream__payload[13:7];
  assign \r_stream__payload.port  = r_stream__payload[17:14];
  assign \r_stream__payload.port.port  = r_stream__payload[16:14];
  assign \r_stream__payload.port.vc_id  = r_stream__payload[17];
  assign \w_stream__payload.new_target  = w_data[13:0];
  assign \w_stream__payload.new_target.target  = w_data[13:0];
  assign \w_stream__payload.new_target.target.x  = w_data[6:0];
  assign \w_stream__payload.new_target.target.y  = w_data[13:7];
  assign \w_stream__payload.port  = w_data[17:14];
  assign \w_stream__payload.port.port  = w_data[16:14];
  assign \w_stream__payload.port.vc_id  = w_data[17];
endmodule

(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:144" *)
(* generator = "Amaranth" *)
module \memory_mapped_router.InputChannel.route_result_fifo.fifo (rst, r_en, w_rdy, r_rdy, r_data, w_en, w_port__data, clk);
  reg \$auto$verilog_backend.cc:2355:dump_module$4  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire [2:0] \$14 ;
  reg \$15 ;
  reg \$16 ;
  reg [1:0] \$17 ;
  wire [1:0] \$2 ;
  wire \$3 ;
  wire [1:0] \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire [2:0] \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* init = 1'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:166" *)
  wire consume;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:141" *)
  reg [1:0] level = 2'h0;
  (* init = 1'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:165" *)
  wire produce;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:241" *)
  output [17:0] r_data;
  wire [17:0] r_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:94" *)
  input r_en;
  wire r_en;
  (* init = 2'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:95" *)
  wire [1:0] r_level;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:240" *)
  reg r_port__addr = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:241" *)
  wire [17:0] r_port__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:93" *)
  output r_rdy;
  wire r_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:87" *)
  wire [17:0] w_data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:89" *)
  input w_en;
  wire w_en;
  (* init = 2'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:90" *)
  wire [1:0] w_level;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:401" *)
  reg w_port__addr = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:87" *)
  input [17:0] w_port__data;
  wire [17:0] w_port__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:400" *)
  wire w_port__en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:88" *)
  output w_rdy;
  wire w_rdy;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:162" *)
  reg [17:0] storage [1:0];
  initial begin
    storage[0] = 18'h00000;
    storage[1] = 18'h00000;
  end
  always @(posedge clk) begin
    if (w_port__en)
      storage[w_port__addr] <= w_port__data;
  end
  assign r_data = storage[r_port__addr];
  assign w_rdy = level != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:153" *) 2'h2;
  assign r_rdy = | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:154" *) level;
  assign w_port__en = w_en & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:171" *) w_rdy;
  assign \$1  = w_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:160" *) w_en;
  assign \$2  = w_port__addr + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:116" *) 1'h1;
  assign \$3  = r_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:159" *) r_en;
  assign \$4  = r_port__addr + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:116" *) 1'h1;
  assign \$5  = w_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:160" *) w_en;
  assign \$6  = r_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:159" *) r_en;
  assign \$7  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:183" *) \$6 ;
  assign \$8  = \$5  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:183" *) \$7 ;
  assign \$9  = level + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:184" *) 1'h1;
  assign \$10  = r_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:159" *) r_en;
  assign \$11  = w_rdy & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:160" *) w_en;
  assign \$12  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:185" *) \$11 ;
  assign \$13  = \$10  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:185" *) \$12 ;
  assign \$14  = level - (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:186" *) 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:165" *)
  always @(posedge clk)
    w_port__addr <= \$15 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:166" *)
  always @(posedge clk)
    r_port__addr <= \$16 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/fifo.py:141" *)
  always @(posedge clk)
    level <= \$17 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$4 ) begin end
    \$15  = w_port__addr;
    if (\$1 ) begin
      \$15  = \$2 [0];
    end
    if (rst) begin
      \$15  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$4 ) begin end
    \$16  = r_port__addr;
    if (\$3 ) begin
      \$16  = \$4 [0];
    end
    if (rst) begin
      \$16  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$4 ) begin end
    \$17  = level;
    if (\$8 ) begin
      \$17  = \$9 [1:0];
    end
    if (\$13 ) begin
      \$17  = \$14 [1:0];
    end
    if (rst) begin
      \$17  = 2'h0;
    end
  end
  assign w_level = level;
  assign r_level = level;
  assign produce = w_port__addr;
  assign w_data = w_port__data;
  assign consume = r_port__addr;
  assign r_port__data = r_data;
endmodule


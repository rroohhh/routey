

package multi_queue_fifo_pkg;

endpackage

interface multi_queue_fifoinput_if import multi_queue_fifo_pkg::*;;
    logic valid;
    logic target;
    logic p;
    logic ready[2];

    modport master (
        output valid,
        output target,
        output p,
        input ready
    );
    modport slave (
        input valid,
        input target,
        input p,
        output ready
    );
    modport monitor (
        input valid,
        input target,
        input p,
        input ready
    );
endinterface

interface multi_queue_fifo_out_stream_if import multi_queue_fifo_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module multi_queue_fifo import multi_queue_fifo_pkg::*;
 (
    input wire clk,
    input wire rst,
    multi_queue_fifoinput_if.slave in,
    multi_queue_fifo_out_stream_if.master out[2]
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueFIFO
    \arq.MultiQueueFIFO  multi_queue_fifo_internal (
        .clk,
        .rst,
        .input__valid(in.valid),
        .input__target(in.target),
        .input__p(in.p),
        .input__ready({<<1{in.ready}}),
        .output__0__payload(out[0].p),
        .output__0__valid(out[0].valid),
        .output__0__ready(out[0].ready),
        .output__1__payload(out[1].p),
        .output__1__valid(out[1].valid),
        .output__1__ready(out[1].ready)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post114, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:636" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueFIFO (input__target, input__p, output__0__ready, output__1__ready, clk, rst, input__ready, output__0__payload, output__0__valid, output__1__payload, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire [4:0] \$1 ;
  wire \$10 ;
  wire [4:0] \$100 ;
  wire \$101 ;
  wire \$102 ;
  wire \$103 ;
  wire [4:0] \$104 ;
  wire \$105 ;
  wire \$106 ;
  wire \$107 ;
  wire \$108 ;
  wire \$109 ;
  wire \$11 ;
  wire \$110 ;
  wire \$111 ;
  wire \$112 ;
  wire \$113 ;
  wire \$114 ;
  wire \$115 ;
  wire \$116 ;
  wire \$117 ;
  wire \$118 ;
  wire \$119 ;
  wire \$12 ;
  wire \$120 ;
  wire \$121 ;
  wire \$122 ;
  wire \$123 ;
  wire \$124 ;
  wire \$125 ;
  wire \$126 ;
  wire \$127 ;
  wire \$128 ;
  wire \$129 ;
  wire \$13 ;
  wire \$130 ;
  wire \$131 ;
  wire \$132 ;
  wire \$133 ;
  wire \$134 ;
  wire \$135 ;
  wire \$136 ;
  wire \$137 ;
  wire \$138 ;
  wire \$139 ;
  wire \$14 ;
  wire \$140 ;
  wire \$141 ;
  wire \$142 ;
  wire \$143 ;
  wire \$144 ;
  wire \$145 ;
  wire [4:0] \$146 ;
  wire \$147 ;
  wire \$148 ;
  wire \$149 ;
  wire \$15 ;
  wire [4:0] \$150 ;
  reg \$151 ;
  reg \$152 ;
  reg \$153 ;
  reg [3:0] \$154 ;
  reg [3:0] \$155 ;
  reg \$156 ;
  reg \$157 ;
  reg \$158 ;
  reg [3:0] \$159 ;
  wire \$16 ;
  reg [3:0] \$160 ;
  wire \$17 ;
  wire \$18 ;
  wire [3:0] \$188 ;
  wire \$19 ;
  wire \$190 ;
  wire [3:0] \$197 ;
  wire \$199 ;
  wire [4:0] \$2 ;
  wire \$20 ;
  wire \$21 ;
  wire \$22 ;
  wire [3:0] \$228 ;
  wire \$23 ;
  wire \$230 ;
  wire [3:0] \$237 ;
  wire \$239 ;
  wire [3:0] \$24 ;
  wire [4:0] \$25 ;
  wire \$26 ;
  wire \$27 ;
  wire \$28 ;
  wire [3:0] \$29 ;
  wire \$3 ;
  wire [4:0] \$30 ;
  wire \$31 ;
  wire \$32 ;
  wire \$33 ;
  wire \$34 ;
  wire \$35 ;
  wire \$36 ;
  wire \$37 ;
  wire \$38 ;
  wire \$39 ;
  wire \$4 ;
  wire \$40 ;
  wire \$41 ;
  wire \$42 ;
  wire \$43 ;
  wire \$44 ;
  wire \$45 ;
  wire \$46 ;
  wire \$47 ;
  wire \$48 ;
  wire \$49 ;
  wire \$5 ;
  wire \$50 ;
  wire \$51 ;
  wire [3:0] \$52 ;
  wire [4:0] \$53 ;
  wire \$54 ;
  wire \$55 ;
  wire \$56 ;
  wire [3:0] \$57 ;
  wire [4:0] \$58 ;
  wire \$59 ;
  wire \$6 ;
  wire \$60 ;
  wire \$61 ;
  wire \$62 ;
  wire \$63 ;
  wire \$64 ;
  wire \$65 ;
  wire \$66 ;
  wire \$67 ;
  wire \$68 ;
  wire \$69 ;
  wire \$7 ;
  wire \$70 ;
  wire \$71 ;
  wire \$72 ;
  wire \$73 ;
  wire \$74 ;
  wire \$75 ;
  wire \$76 ;
  wire \$77 ;
  wire \$78 ;
  wire \$79 ;
  wire \$8 ;
  wire \$80 ;
  wire \$81 ;
  wire \$82 ;
  wire \$83 ;
  wire \$84 ;
  wire \$85 ;
  wire \$86 ;
  wire \$87 ;
  wire \$88 ;
  wire \$89 ;
  wire \$9 ;
  wire \$90 ;
  wire \$91 ;
  wire \$92 ;
  wire \$93 ;
  wire \$94 ;
  wire \$95 ;
  wire \$96 ;
  wire \$97 ;
  wire \$98 ;
  wire \$99 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:236" *)
  reg [3:0] buffer_read__addr;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:237" *)
  wire buffer_read__data;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:235" *)
  reg buffer_read__en;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:397" *)
  reg [3:0] buffer_write__addr;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:398" *)
  reg buffer_write__data;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:396" *)
  reg buffer_write__en;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:607" *)
  input input__p;
  wire input__p;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:625" *)
  output [1:0] input__ready;
  wire [1:0] input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:625" *)
  wire \input__ready[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:625" *)
  wire \input__ready[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:606" *)
  input input__target;
  wire input__target;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:605" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:657" *)
  reg mem_out_have_data = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:658" *)
  reg mem_out_id = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:640" *)
  reg out_reg_0 = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:640" *)
  reg out_reg_1 = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:641" *)
  reg out_reg_filled_0 = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:641" *)
  reg out_reg_filled_1 = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__0__payload;
  wire output__0__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__1__payload;
  wire output__1__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* capacity = 32'd8 *)
  (* debug_item = 32'd1 *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:643" *)
  wire [3:0] outstanding_0;
  (* capacity = 32'd8 *)
  (* debug_item = 32'd1 *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:643" *)
  wire [3:0] outstanding_1;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:686" *)
  wire pop_0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:686" *)
  wire pop_1;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:684" *)
  wire push_0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:684" *)
  wire push_1;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:638" *)
  reg [3:0] read_ptr_0 = 4'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:638" *)
  reg [3:0] read_ptr_1 = 4'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:639" *)
  reg [3:0] write_ptr_0 = 4'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:639" *)
  reg [3:0] write_ptr_1 = 4'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:650" *)
  reg [0:0] buffer [15:0];
  initial begin
    buffer[0] = 1'h0;
    buffer[1] = 1'h0;
    buffer[2] = 1'h0;
    buffer[3] = 1'h0;
    buffer[4] = 1'h0;
    buffer[5] = 1'h0;
    buffer[6] = 1'h0;
    buffer[7] = 1'h0;
    buffer[8] = 1'h0;
    buffer[9] = 1'h0;
    buffer[10] = 1'h0;
    buffer[11] = 1'h0;
    buffer[12] = 1'h0;
    buffer[13] = 1'h0;
    buffer[14] = 1'h0;
    buffer[15] = 1'h0;
  end
  always @(posedge clk) begin
    if (buffer_write__en)
      buffer[buffer_write__addr] <= buffer_write__data;
  end
  reg [0:0] _0_;
  always @(posedge clk) begin
    if (buffer_read__en) begin
      _0_ <= buffer[buffer_read__addr];
    end
  end
  assign buffer_read__data = _0_;
  assign \$1  = write_ptr_0 - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:645" *) read_ptr_0;
  assign \$2  = write_ptr_1 - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:645" *) read_ptr_1;
  assign \$3  = input__ready[0] & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:685" *) input__valid;
  assign \$4  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:685" *) input__target;
  assign push_0 = \$3  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:685" *) \$4 ;
  assign pop_0 = output__0__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:687" *) output__0__valid;
  assign \$5  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) mem_out_id;
  assign \$6  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$5 ;
  assign output__0__valid = out_reg_filled_0 | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:724" *) \$6 ;
  assign output__0__payload = out_reg_filled_0 ? (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:725" *) out_reg_0 : buffer_read__data;
  assign \$7  = read_ptr_0[3] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:682" *) write_ptr_0[3];
  assign \$8  = read_ptr_0[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:682" *) write_ptr_0[2:0];
  assign \$9  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:682" *) \$8 ;
  assign \$10  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:726" *) \$9 ;
  assign \$11  = read_ptr_0 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_0;
  assign \$12  = push_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$11 ;
  assign \$13  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_0;
  assign \$14  = \$13  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$15  = \$12  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$14 ;
  assign \$16  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) mem_out_id;
  assign \$17  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$16 ;
  assign \$18  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$19  = \$17  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$18 ;
  assign \$20  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$19 ;
  assign \$21  = \$15  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$20 ;
  assign \$22  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$21 ;
  assign \$23  = push_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$22 ;
  assign \$188  = write_ptr_0 % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:733" *) 4'h8;
  assign \$25  = 1'h0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:733" *) \$24 ;
  assign \$26  = read_ptr_0 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_0;
  assign \$27  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$26 ;
  assign \$28  = pop_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$27 ;
  assign \$197  = read_ptr_0 % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:667" *) 4'h8;
  assign \$30  = 1'h0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:667" *) \$29 ;
  assign \$31  = input__ready[1] & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:685" *) input__valid;
  assign push_1 = \$31  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:685" *) \$32 ;
  assign pop_1 = output__1__ready & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:687" *) output__1__valid;
  assign \$34  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$33 ;
  assign output__1__valid = out_reg_filled_1 | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:724" *) \$34 ;
  assign output__1__payload = out_reg_filled_1 ? (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:725" *) out_reg_1 : buffer_read__data;
  assign \$35  = read_ptr_1[3] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:682" *) write_ptr_1[3];
  assign \$36  = read_ptr_1[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:682" *) write_ptr_1[2:0];
  assign \$37  = \$35  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:682" *) \$36 ;
  assign \$38  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:726" *) \$37 ;
  assign \$39  = read_ptr_1 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_1;
  assign \$40  = push_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$39 ;
  assign \$41  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_1;
  assign \$42  = \$41  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$43  = \$40  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$42 ;
  assign \$45  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$44 ;
  assign \$46  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$47  = \$45  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$46 ;
  assign \$48  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$47 ;
  assign \$49  = \$43  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$48 ;
  assign \$50  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$49 ;
  assign \$51  = push_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$50 ;
  assign \$228  = write_ptr_1 % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:733" *) 4'h8;
  assign \$53  = 4'h8 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:733" *) \$52 ;
  assign \$54  = read_ptr_1 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_1;
  assign \$55  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$54 ;
  assign \$56  = pop_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$55 ;
  assign \$237  = read_ptr_1 % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:667" *) 4'h8;
  assign \$58  = 4'h8 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:667" *) \$57 ;
  assign \$59  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) mem_out_id;
  assign \$60  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$59 ;
  assign \$61  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:703" *) pop_0;
  assign \$62  = \$60  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:703" *) \$61 ;
  assign \$63  = read_ptr_0 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_0;
  assign \$64  = push_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$63 ;
  assign \$65  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_0;
  assign \$66  = \$65  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$67  = \$64  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$66 ;
  assign \$68  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) mem_out_id;
  assign \$69  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$68 ;
  assign \$70  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$71  = \$69  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$70 ;
  assign \$72  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$71 ;
  assign \$73  = \$67  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$72 ;
  assign \$74  = read_ptr_0 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_0;
  assign \$75  = push_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$74 ;
  assign \$76  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_0;
  assign \$77  = \$76  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$78  = \$75  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$77 ;
  assign \$79  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) mem_out_id;
  assign \$80  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$79 ;
  assign \$81  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$82  = \$80  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$81 ;
  assign \$83  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$82 ;
  assign \$84  = \$78  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$83 ;
  assign \$85  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:717" *) \$84 ;
  assign \$86  = pop_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:717" *) \$85 ;
  assign \$87  = read_ptr_0 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_0;
  assign \$88  = push_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$87 ;
  assign \$89  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_0;
  assign \$90  = \$89  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$91  = \$88  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$90 ;
  assign \$92  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) mem_out_id;
  assign \$93  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$92 ;
  assign \$94  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_0;
  assign \$95  = \$93  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$94 ;
  assign \$96  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$95 ;
  assign \$97  = \$91  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$96 ;
  assign \$98  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$97 ;
  assign \$99  = push_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$98 ;
  assign \$100  = write_ptr_0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:673" *) 1'h1;
  assign \$101  = read_ptr_0 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_0;
  assign \$102  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$101 ;
  assign \$103  = pop_0 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$102 ;
  assign \$104  = read_ptr_0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:673" *) 1'h1;
  assign \$106  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$105 ;
  assign \$107  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:703" *) pop_1;
  assign \$108  = \$106  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:703" *) \$107 ;
  assign \$109  = read_ptr_1 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_1;
  assign \$110  = push_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$109 ;
  assign \$111  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_1;
  assign \$112  = \$111  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$113  = \$110  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$112 ;
  assign \$115  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$114 ;
  assign \$116  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$117  = \$115  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$116 ;
  assign \$118  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$117 ;
  assign \$119  = \$113  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$118 ;
  assign \$120  = read_ptr_1 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_1;
  assign \$121  = push_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$120 ;
  assign \$122  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_1;
  assign \$123  = \$122  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$124  = \$121  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$123 ;
  assign \$126  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$125 ;
  assign \$127  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$128  = \$126  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$127 ;
  assign \$129  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$128 ;
  assign \$130  = \$124  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$129 ;
  assign \$131  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:717" *) \$130 ;
  assign \$132  = pop_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:717" *) \$131 ;
  assign \$133  = read_ptr_1 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_1;
  assign \$134  = push_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$133 ;
  assign \$135  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) out_reg_filled_1;
  assign \$136  = \$135  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$137  = \$134  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$136 ;
  assign \$139  = mem_out_have_data & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:689" *) \$138 ;
  assign \$140  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) pop_1;
  assign \$141  = \$139  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$140 ;
  assign \$142  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$141 ;
  assign \$143  = \$137  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:696" *) \$142 ;
  assign \$144  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$143 ;
  assign \$145  = push_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:697" *) \$144 ;
  assign \$146  = write_ptr_1 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:673" *) 1'h1;
  assign \$147  = read_ptr_1 == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:681" *) write_ptr_1;
  assign \$148  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$147 ;
  assign \$149  = pop_1 & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:700" *) \$148 ;
  assign \$150  = read_ptr_1 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:673" *) 1'h1;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:657" *)
  always @(posedge clk)
    mem_out_have_data <= \$151 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:641" *)
  always @(posedge clk)
    out_reg_filled_0 <= \$152 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:640" *)
  always @(posedge clk)
    out_reg_0 <= \$153 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:639" *)
  always @(posedge clk)
    write_ptr_0 <= \$154 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:638" *)
  always @(posedge clk)
    read_ptr_0 <= \$155 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:658" *)
  always @(posedge clk)
    mem_out_id <= \$156 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:641" *)
  always @(posedge clk)
    out_reg_filled_1 <= \$157 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:640" *)
  always @(posedge clk)
    out_reg_1 <= \$158 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:639" *)
  always @(posedge clk)
    write_ptr_1 <= \$159 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:638" *)
  always @(posedge clk)
    read_ptr_1 <= \$160 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_read__en = 1'h0;
    if (\$28 ) begin
      buffer_read__en = 1'h1;
    end
    if (\$56 ) begin
      buffer_read__en = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_write__addr = 4'h0;
    if (\$23 ) begin
      buffer_write__addr = \$25 [3:0];
    end
    if (\$51 ) begin
      buffer_write__addr = \$53 [3:0];
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_write__en = 1'h0;
    if (\$23 ) begin
      buffer_write__en = 1'h1;
    end
    if (\$51 ) begin
      buffer_write__en = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_write__data = 1'h0;
    if (\$23 ) begin
      buffer_write__data = input__p;
    end
    if (\$51 ) begin
      buffer_write__data = input__p;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_read__addr = 4'h0;
    if (\$28 ) begin
      buffer_read__addr = \$30 [3:0];
    end
    if (\$56 ) begin
      buffer_read__addr = \$58 [3:0];
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$151  = buffer_read__en;
    if (rst) begin
      \$151  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$152  = out_reg_filled_0;
    if (\$62 ) begin
      \$152  = 1'h1;
    end
    if (\$73 ) begin
      \$152  = 1'h1;
    end
    if (\$86 ) begin
      \$152  = 1'h0;
    end
    if (rst) begin
      \$152  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$153  = out_reg_0;
    if (\$62 ) begin
      \$153  = buffer_read__data;
    end
    if (\$73 ) begin
      \$153  = input__p;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$154  = write_ptr_0;
    if (\$99 ) begin
      \$154  = \$100 [3:0];
    end
    if (rst) begin
      \$154  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$155  = read_ptr_0;
    if (\$103 ) begin
      \$155  = \$104 [3:0];
    end
    if (rst) begin
      \$155  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$156  = mem_out_id;
    if (\$103 ) begin
      \$156  = 1'h0;
    end
    if (\$149 ) begin
      \$156  = 1'h1;
    end
    if (rst) begin
      \$156  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$157  = out_reg_filled_1;
    if (\$108 ) begin
      \$157  = 1'h1;
    end
    if (\$119 ) begin
      \$157  = 1'h1;
    end
    if (\$132 ) begin
      \$157  = 1'h0;
    end
    if (rst) begin
      \$157  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$158  = out_reg_1;
    if (\$108 ) begin
      \$158  = buffer_read__data;
    end
    if (\$119 ) begin
      \$158  = input__p;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$159  = write_ptr_1;
    if (\$145 ) begin
      \$159  = \$146 [3:0];
    end
    if (rst) begin
      \$159  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$160  = read_ptr_1;
    if (\$149 ) begin
      \$160  = \$150 [3:0];
    end
    if (rst) begin
      \$160  = 4'h0;
    end
  end
  assign outstanding_0 = \$1 [3:0];
  assign outstanding_1 = \$2 [3:0];
  assign \input__ready[0]  = input__ready[0];
  assign \input__ready[1]  = input__ready[1];
  assign input__ready[1] = \$38 ;
  assign input__ready[0] = \$10 ;
  assign \$190  = 1'h1;
  assign \$24  = \$188 ;
  assign \$199  = 1'h1;
  assign \$29  = \$197 ;
  assign \$32  = input__target;
  assign \$33  = mem_out_id;
  assign \$44  = mem_out_id;
  assign \$230  = 1'h1;
  assign \$52  = \$228 ;
  assign \$239  = 1'h1;
  assign \$57  = \$237 ;
  assign \$105  = mem_out_id;
  assign \$114  = mem_out_id;
  assign \$125  = mem_out_id;
  assign \$138  = mem_out_id;
endmodule


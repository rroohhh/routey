

package multi_queue_credit_counter_rx_pkg;
typedef struct packed {
    logic ready;
    logic valid;
} stream_monitor;
endpackage

interface multi_queue_credit_counter_rx_credit_out_if import multi_queue_credit_counter_rx_pkg::*;;
    logic [3: 0] credit[2];
    logic did_trigger;
    logic trigger;

    modport master (
        output credit,
        input did_trigger,
        output trigger
    );
    modport slave (
        input credit,
        output did_trigger,
        input trigger
    );
    modport monitor (
        input credit,
        input did_trigger,
        input trigger
    );
endinterface

module multi_queue_credit_counter_rx import multi_queue_credit_counter_rx_pkg::*;
 (
    input wire clk,
    input wire rst,
    input wire stream_monitor fifo_output_monitor[2],
    multi_queue_credit_counter_rx_credit_out_if.master credit_out
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueCreditCounterRX
    \arq.MultiQueueCreditCounterRX  multi_queue_credit_counter_rx_internal (
        .clk,
        .rst,
        .fifo_output_monitor__0(fifo_output_monitor[0]),
        .fifo_output_monitor__1(fifo_output_monitor[1]),
        .credit_out__credit({<<4{credit_out.credit}}),
        .credit_out__did_trigger(credit_out.did_trigger),
        .credit_out__trigger(credit_out.trigger)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:839" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueCreditCounterRX (fifo_output_monitor__1, credit_out__did_trigger, clk, rst, credit_out__credit, credit_out__trigger, fifo_output_monitor__0);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  reg \$10 ;
  wire \$2 ;
  wire [4:0] \$3 ;
  wire \$4 ;
  wire [4:0] \$5 ;
  wire \$6 ;
  wire [1:0] \$7 ;
  reg [3:0] \$8 ;
  reg [3:0] \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:830" *)
  output [7:0] credit_out__credit;
  wire [7:0] credit_out__credit;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:830" *)
  wire [3:0] \credit_out__credit[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:830" *)
  wire [3:0] \credit_out__credit[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:823" *)
  input credit_out__did_trigger;
  wire credit_out__did_trigger;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:824" *)
  output credit_out__trigger;
  reg credit_out__trigger;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:849" *)
  reg credit_trigger_timer = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  input [1:0] fifo_output_monitor__0;
  wire [1:0] fifo_output_monitor__0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__0.ready ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__0.valid ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  input [1:0] fifo_output_monitor__1;
  wire [1:0] fifo_output_monitor__1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__1.ready ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__1.valid ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:841" *)
  reg [3:0] read_ptr_0 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:841" *)
  reg [3:0] read_ptr_1 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  assign \$2  = fifo_output_monitor__0[0] & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:845" *) fifo_output_monitor__0[1];
  assign \$3  = read_ptr_0 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:846" *) 1'h1;
  assign \$4  = fifo_output_monitor__1[0] & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:845" *) fifo_output_monitor__1[1];
  assign \$5  = read_ptr_1 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:846" *) 1'h1;
  assign \$7  = credit_trigger_timer + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:858" *) 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:841" *)
  always @(posedge clk)
    read_ptr_0 <= \$8 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:841" *)
  always @(posedge clk)
    read_ptr_1 <= \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:849" *)
  always @(posedge clk)
    credit_trigger_timer <= \$10 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    credit_out__trigger = 1'h0;
    (* full_case = 32'd1 *)
    if (credit_out__did_trigger) begin
    end else begin
      if (\$1 ) begin
        credit_out__trigger = 1'h1;
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$8  = read_ptr_0;
    if (\$2 ) begin
      \$8  = \$3 [3:0];
    end
    if (rst) begin
      \$8  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$9  = read_ptr_1;
    if (\$4 ) begin
      \$9  = \$5 [3:0];
    end
    if (rst) begin
      \$9  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (credit_out__did_trigger) begin
      \$10  = 1'h0;
    end else begin
      (* full_case = 32'd1 *)
      if (\$6 ) begin
        \$10  = 1'h0;
      end else begin
        \$10  = \$7 [0];
      end
    end
    if (rst) begin
      \$10  = 1'h0;
    end
  end
  assign \fifo_output_monitor__0.valid  = fifo_output_monitor__0[0];
  assign \fifo_output_monitor__0.ready  = fifo_output_monitor__0[1];
  assign \fifo_output_monitor__1.valid  = fifo_output_monitor__1[0];
  assign \fifo_output_monitor__1.ready  = fifo_output_monitor__1[1];
  assign \credit_out__credit[0]  = credit_out__credit[3:0];
  assign \credit_out__credit[1]  = credit_out__credit[7:4];
  assign credit_out__credit[7:4] = read_ptr_1;
  assign credit_out__credit[3:0] = read_ptr_0;
  assign \$1  = credit_trigger_timer;
  assign \$6  = credit_trigger_timer;
endmodule




package multi_queue_fifo_pkg;

endpackage

interface multi_queue_fifo_in_if import multi_queue_fifo_pkg::*;;
    logic valid;
    logic target;
    logic p;
    logic ready[2];

    modport master (
        output valid,
        output target,
        output p,
        input ready
    );
    modport slave (
        input valid,
        input target,
        input p,
        output ready
    );
    modport monitor (
        input valid,
        input target,
        input p,
        input ready
    );
endinterface

interface multi_queue_fifo_out_stream_if import multi_queue_fifo_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module multi_queue_fifo import multi_queue_fifo_pkg::*;
 (
    input wire clk,
    input wire rst,
    multi_queue_fifo_in_if.slave in,
    multi_queue_fifo_out_stream_if.master out[2]
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueFIFO
    \arq.MultiQueueFIFO  multi_queue_fifo_internal (
        .clk,
        .rst,
        .input__valid(in.valid),
        .input__target(in.target),
        .input__p(in.p),
        .input__ready({<<1{in.ready}}),
        .output__0__payload(out[0].p),
        .output__0__valid(out[0].valid),
        .output__0__ready(out[0].ready),
        .output__1__payload(out[1].p),
        .output__1__valid(out[1].valid),
        .output__1__ready(out[1].ready)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:558" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueFIFO (input__target, input__p, output__0__ready, output__1__ready, clk, rst, input__ready, output__0__payload, output__0__valid, output__1__payload, output__1__valid, input__valid);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$100 ;
  wire \$101 ;
  wire [4:0] \$102 ;
  wire \$103 ;
  wire \$104 ;
  wire \$105 ;
  wire \$106 ;
  wire \$107 ;
  wire \$108 ;
  wire \$109 ;
  wire \$11 ;
  wire \$110 ;
  wire \$111 ;
  wire \$112 ;
  wire \$113 ;
  wire \$114 ;
  wire \$115 ;
  wire \$116 ;
  wire \$117 ;
  wire \$118 ;
  wire \$119 ;
  wire \$12 ;
  wire \$120 ;
  wire \$121 ;
  wire \$122 ;
  wire \$123 ;
  wire \$124 ;
  wire \$125 ;
  wire \$126 ;
  wire \$127 ;
  wire \$128 ;
  wire \$129 ;
  wire \$13 ;
  wire \$130 ;
  wire \$131 ;
  wire \$132 ;
  wire \$133 ;
  wire \$134 ;
  wire \$135 ;
  wire \$136 ;
  wire \$137 ;
  wire \$138 ;
  wire \$139 ;
  wire \$14 ;
  wire \$140 ;
  wire \$141 ;
  wire \$142 ;
  wire \$143 ;
  wire [4:0] \$144 ;
  wire \$145 ;
  wire \$146 ;
  wire \$147 ;
  wire [4:0] \$148 ;
  reg \$149 ;
  wire \$15 ;
  reg \$150 ;
  reg \$151 ;
  reg [3:0] \$152 ;
  reg [3:0] \$153 ;
  reg \$154 ;
  reg \$155 ;
  reg \$156 ;
  reg [3:0] \$157 ;
  reg [3:0] \$158 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire [3:0] \$184 ;
  wire \$186 ;
  wire \$19 ;
  wire [3:0] \$193 ;
  wire \$195 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  wire [3:0] \$22 ;
  wire [3:0] \$224 ;
  wire \$226 ;
  wire [4:0] \$23 ;
  wire [3:0] \$233 ;
  wire \$235 ;
  wire \$24 ;
  wire \$25 ;
  wire \$26 ;
  wire [3:0] \$27 ;
  wire [4:0] \$28 ;
  wire \$29 ;
  wire \$3 ;
  wire \$30 ;
  wire \$31 ;
  wire \$32 ;
  wire \$33 ;
  wire \$34 ;
  wire \$35 ;
  wire \$36 ;
  wire \$37 ;
  wire \$38 ;
  wire \$39 ;
  wire \$4 ;
  wire \$40 ;
  wire \$41 ;
  wire \$42 ;
  wire \$43 ;
  wire \$44 ;
  wire \$45 ;
  wire \$46 ;
  wire \$47 ;
  wire \$48 ;
  wire \$49 ;
  wire \$5 ;
  wire [3:0] \$50 ;
  wire [4:0] \$51 ;
  wire \$52 ;
  wire \$53 ;
  wire \$54 ;
  wire [3:0] \$55 ;
  wire [4:0] \$56 ;
  wire \$57 ;
  wire \$58 ;
  wire \$59 ;
  wire \$6 ;
  wire \$60 ;
  wire \$61 ;
  wire \$62 ;
  wire \$63 ;
  wire \$64 ;
  wire \$65 ;
  wire \$66 ;
  wire \$67 ;
  wire \$68 ;
  wire \$69 ;
  wire \$7 ;
  wire \$70 ;
  wire \$71 ;
  wire \$72 ;
  wire \$73 ;
  wire \$74 ;
  wire \$75 ;
  wire \$76 ;
  wire \$77 ;
  wire \$78 ;
  wire \$79 ;
  wire \$8 ;
  wire \$80 ;
  wire \$81 ;
  wire \$82 ;
  wire \$83 ;
  wire \$84 ;
  wire \$85 ;
  wire \$86 ;
  wire \$87 ;
  wire \$88 ;
  wire \$89 ;
  wire \$9 ;
  wire \$90 ;
  wire \$91 ;
  wire \$92 ;
  wire \$93 ;
  wire \$94 ;
  wire \$95 ;
  wire \$96 ;
  wire \$97 ;
  wire [4:0] \$98 ;
  wire \$99 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:240" *)
  reg [3:0] buffer_read__addr;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:241" *)
  wire buffer_read__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:239" *)
  reg buffer_read__en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:401" *)
  reg [3:0] buffer_write__addr;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:402" *)
  reg buffer_write__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:400" *)
  reg buffer_write__en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:538" *)
  input input__p;
  wire input__p;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:547" *)
  output [1:0] input__ready;
  wire [1:0] input__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:547" *)
  wire \input__ready[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:547" *)
  wire \input__ready[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:537" *)
  input input__target;
  wire input__target;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:536" *)
  input input__valid;
  wire input__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:572" *)
  reg mem_out_have_data = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:573" *)
  reg mem_out_id = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:562" *)
  reg out_reg_0 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:562" *)
  reg out_reg_1 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:563" *)
  reg out_reg_filled_0 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:563" *)
  reg out_reg_filled_1 = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__0__payload;
  wire output__0__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__0__ready;
  wire output__0__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__0__valid;
  wire output__0__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__1__payload;
  wire output__1__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__1__ready;
  wire output__1__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__1__valid;
  wire output__1__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:601" *)
  wire pop_0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:601" *)
  wire pop_1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:599" *)
  wire push_0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:599" *)
  wire push_1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:560" *)
  reg [3:0] read_ptr_0 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:560" *)
  reg [3:0] read_ptr_1 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:561" *)
  reg [3:0] write_ptr_0 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:561" *)
  reg [3:0] write_ptr_1 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:565" *)
  reg [0:0] buffer [15:0];
  initial begin
    buffer[0] = 1'h0;
    buffer[1] = 1'h0;
    buffer[2] = 1'h0;
    buffer[3] = 1'h0;
    buffer[4] = 1'h0;
    buffer[5] = 1'h0;
    buffer[6] = 1'h0;
    buffer[7] = 1'h0;
    buffer[8] = 1'h0;
    buffer[9] = 1'h0;
    buffer[10] = 1'h0;
    buffer[11] = 1'h0;
    buffer[12] = 1'h0;
    buffer[13] = 1'h0;
    buffer[14] = 1'h0;
    buffer[15] = 1'h0;
  end
  always @(posedge clk) begin
    if (buffer_write__en)
      buffer[buffer_write__addr] <= buffer_write__data;
  end
  reg [0:0] _0_;
  always @(posedge clk) begin
    if (buffer_read__en) begin
      _0_ <= buffer[buffer_read__addr];
    end
  end
  assign buffer_read__data = _0_;
  assign \$1  = input__ready[0] & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:600" *) input__valid;
  assign \$2  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:600" *) input__target;
  assign push_0 = \$1  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:600" *) \$2 ;
  assign pop_0 = output__0__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:602" *) output__0__valid;
  assign \$3  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) mem_out_id;
  assign \$4  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$3 ;
  assign output__0__valid = out_reg_filled_0 | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:639" *) \$4 ;
  assign output__0__payload = out_reg_filled_0 ? (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:640" *) out_reg_0 : buffer_read__data;
  assign \$5  = read_ptr_0[3] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:597" *) write_ptr_0[3];
  assign \$6  = read_ptr_0[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:597" *) write_ptr_0[2:0];
  assign \$7  = \$5  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:597" *) \$6 ;
  assign \$8  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:641" *) \$7 ;
  assign \$9  = read_ptr_0 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_0;
  assign \$10  = push_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$9 ;
  assign \$11  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_0;
  assign \$12  = \$11  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$13  = \$10  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$12 ;
  assign \$14  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) mem_out_id;
  assign \$15  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$14 ;
  assign \$16  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$17  = \$15  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$16 ;
  assign \$18  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$17 ;
  assign \$19  = \$13  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$18 ;
  assign \$20  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$19 ;
  assign \$21  = push_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$20 ;
  assign \$184  = write_ptr_0 % (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:648" *) 4'h8;
  assign \$23  = 1'h0 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:648" *) \$22 ;
  assign \$24  = read_ptr_0 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_0;
  assign \$25  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$24 ;
  assign \$26  = pop_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$25 ;
  assign \$193  = read_ptr_0 % (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:582" *) 4'h8;
  assign \$28  = 1'h0 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:582" *) \$27 ;
  assign \$29  = input__ready[1] & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:600" *) input__valid;
  assign push_1 = \$29  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:600" *) \$30 ;
  assign pop_1 = output__1__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:602" *) output__1__valid;
  assign \$32  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$31 ;
  assign output__1__valid = out_reg_filled_1 | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:639" *) \$32 ;
  assign output__1__payload = out_reg_filled_1 ? (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:640" *) out_reg_1 : buffer_read__data;
  assign \$33  = read_ptr_1[3] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:597" *) write_ptr_1[3];
  assign \$34  = read_ptr_1[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:597" *) write_ptr_1[2:0];
  assign \$35  = \$33  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:597" *) \$34 ;
  assign \$36  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:641" *) \$35 ;
  assign \$37  = read_ptr_1 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_1;
  assign \$38  = push_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$37 ;
  assign \$39  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_1;
  assign \$40  = \$39  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$41  = \$38  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$40 ;
  assign \$43  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$42 ;
  assign \$44  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$45  = \$43  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$44 ;
  assign \$46  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$45 ;
  assign \$47  = \$41  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$46 ;
  assign \$48  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$47 ;
  assign \$49  = push_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$48 ;
  assign \$224  = write_ptr_1 % (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:648" *) 4'h8;
  assign \$51  = 4'h8 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:648" *) \$50 ;
  assign \$52  = read_ptr_1 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_1;
  assign \$53  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$52 ;
  assign \$54  = pop_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$53 ;
  assign \$233  = read_ptr_1 % (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:582" *) 4'h8;
  assign \$56  = 4'h8 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:582" *) \$55 ;
  assign \$57  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) mem_out_id;
  assign \$58  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$57 ;
  assign \$59  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:618" *) pop_0;
  assign \$60  = \$58  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:618" *) \$59 ;
  assign \$61  = read_ptr_0 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_0;
  assign \$62  = push_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$61 ;
  assign \$63  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_0;
  assign \$64  = \$63  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$65  = \$62  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$64 ;
  assign \$66  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) mem_out_id;
  assign \$67  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$66 ;
  assign \$68  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$69  = \$67  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$68 ;
  assign \$70  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$69 ;
  assign \$71  = \$65  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$70 ;
  assign \$72  = read_ptr_0 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_0;
  assign \$73  = push_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$72 ;
  assign \$74  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_0;
  assign \$75  = \$74  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$76  = \$73  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$75 ;
  assign \$77  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) mem_out_id;
  assign \$78  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$77 ;
  assign \$79  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$80  = \$78  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$79 ;
  assign \$81  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$80 ;
  assign \$82  = \$76  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$81 ;
  assign \$83  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:632" *) \$82 ;
  assign \$84  = pop_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:632" *) \$83 ;
  assign \$85  = read_ptr_0 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_0;
  assign \$86  = push_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$85 ;
  assign \$87  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_0;
  assign \$88  = \$87  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$89  = \$86  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$88 ;
  assign \$90  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) mem_out_id;
  assign \$91  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$90 ;
  assign \$92  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_0;
  assign \$93  = \$91  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$92 ;
  assign \$94  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$93 ;
  assign \$95  = \$89  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$94 ;
  assign \$96  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$95 ;
  assign \$97  = push_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$96 ;
  assign \$98  = write_ptr_0 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:588" *) 1'h1;
  assign \$99  = read_ptr_0 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_0;
  assign \$100  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$99 ;
  assign \$101  = pop_0 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$100 ;
  assign \$102  = read_ptr_0 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:588" *) 1'h1;
  assign \$104  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$103 ;
  assign \$105  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:618" *) pop_1;
  assign \$106  = \$104  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:618" *) \$105 ;
  assign \$107  = read_ptr_1 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_1;
  assign \$108  = push_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$107 ;
  assign \$109  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_1;
  assign \$110  = \$109  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$111  = \$108  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$110 ;
  assign \$113  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$112 ;
  assign \$114  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$115  = \$113  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$114 ;
  assign \$116  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$115 ;
  assign \$117  = \$111  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$116 ;
  assign \$118  = read_ptr_1 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_1;
  assign \$119  = push_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$118 ;
  assign \$120  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_1;
  assign \$121  = \$120  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$122  = \$119  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$121 ;
  assign \$124  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$123 ;
  assign \$125  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$126  = \$124  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$125 ;
  assign \$127  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$126 ;
  assign \$128  = \$122  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$127 ;
  assign \$129  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:632" *) \$128 ;
  assign \$130  = pop_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:632" *) \$129 ;
  assign \$131  = read_ptr_1 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_1;
  assign \$132  = push_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$131 ;
  assign \$133  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) out_reg_filled_1;
  assign \$134  = \$133  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$135  = \$132  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$134 ;
  assign \$137  = mem_out_have_data & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:604" *) \$136 ;
  assign \$138  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) pop_1;
  assign \$139  = \$137  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$138 ;
  assign \$140  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$139 ;
  assign \$141  = \$135  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:611" *) \$140 ;
  assign \$142  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$141 ;
  assign \$143  = push_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:612" *) \$142 ;
  assign \$144  = write_ptr_1 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:588" *) 1'h1;
  assign \$145  = read_ptr_1 == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:596" *) write_ptr_1;
  assign \$146  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$145 ;
  assign \$147  = pop_1 & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:615" *) \$146 ;
  assign \$148  = read_ptr_1 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:588" *) 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:572" *)
  always @(posedge clk)
    mem_out_have_data <= \$149 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:563" *)
  always @(posedge clk)
    out_reg_filled_0 <= \$150 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:562" *)
  always @(posedge clk)
    out_reg_0 <= \$151 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:561" *)
  always @(posedge clk)
    write_ptr_0 <= \$152 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:560" *)
  always @(posedge clk)
    read_ptr_0 <= \$153 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:573" *)
  always @(posedge clk)
    mem_out_id <= \$154 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:563" *)
  always @(posedge clk)
    out_reg_filled_1 <= \$155 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:562" *)
  always @(posedge clk)
    out_reg_1 <= \$156 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:561" *)
  always @(posedge clk)
    write_ptr_1 <= \$157 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:560" *)
  always @(posedge clk)
    read_ptr_1 <= \$158 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_read__en = 1'h0;
    if (\$26 ) begin
      buffer_read__en = 1'h1;
    end
    if (\$54 ) begin
      buffer_read__en = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_write__addr = 4'h0;
    if (\$21 ) begin
      buffer_write__addr = \$23 [3:0];
    end
    if (\$49 ) begin
      buffer_write__addr = \$51 [3:0];
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_write__en = 1'h0;
    if (\$21 ) begin
      buffer_write__en = 1'h1;
    end
    if (\$49 ) begin
      buffer_write__en = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_write__data = 1'h0;
    if (\$21 ) begin
      buffer_write__data = input__p;
    end
    if (\$49 ) begin
      buffer_write__data = input__p;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    buffer_read__addr = 4'h0;
    if (\$26 ) begin
      buffer_read__addr = \$28 [3:0];
    end
    if (\$54 ) begin
      buffer_read__addr = \$56 [3:0];
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$149  = buffer_read__en;
    if (rst) begin
      \$149  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$150  = out_reg_filled_0;
    if (\$60 ) begin
      \$150  = 1'h1;
    end
    if (\$71 ) begin
      \$150  = 1'h1;
    end
    if (\$84 ) begin
      \$150  = 1'h0;
    end
    if (rst) begin
      \$150  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$151  = out_reg_0;
    if (\$60 ) begin
      \$151  = buffer_read__data;
    end
    if (\$71 ) begin
      \$151  = input__p;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$152  = write_ptr_0;
    if (\$97 ) begin
      \$152  = \$98 [3:0];
    end
    if (rst) begin
      \$152  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$153  = read_ptr_0;
    if (\$101 ) begin
      \$153  = \$102 [3:0];
    end
    if (rst) begin
      \$153  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$154  = mem_out_id;
    if (\$101 ) begin
      \$154  = 1'h0;
    end
    if (\$147 ) begin
      \$154  = 1'h1;
    end
    if (rst) begin
      \$154  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$155  = out_reg_filled_1;
    if (\$106 ) begin
      \$155  = 1'h1;
    end
    if (\$117 ) begin
      \$155  = 1'h1;
    end
    if (\$130 ) begin
      \$155  = 1'h0;
    end
    if (rst) begin
      \$155  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$156  = out_reg_1;
    if (\$106 ) begin
      \$156  = buffer_read__data;
    end
    if (\$117 ) begin
      \$156  = input__p;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$157  = write_ptr_1;
    if (\$143 ) begin
      \$157  = \$144 [3:0];
    end
    if (rst) begin
      \$157  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$158  = read_ptr_1;
    if (\$147 ) begin
      \$158  = \$148 [3:0];
    end
    if (rst) begin
      \$158  = 4'h0;
    end
  end
  assign \input__ready[0]  = input__ready[0];
  assign \input__ready[1]  = input__ready[1];
  assign input__ready[1] = \$36 ;
  assign input__ready[0] = \$8 ;
  assign \$186  = 1'h1;
  assign \$22  = \$184 ;
  assign \$195  = 1'h1;
  assign \$27  = \$193 ;
  assign \$30  = input__target;
  assign \$31  = mem_out_id;
  assign \$42  = mem_out_id;
  assign \$226  = 1'h1;
  assign \$50  = \$224 ;
  assign \$235  = 1'h1;
  assign \$55  = \$233 ;
  assign \$103  = mem_out_id;
  assign \$112  = mem_out_id;
  assign \$123  = mem_out_id;
  assign \$136  = mem_out_id;
endmodule




package lwwreg_pkg;

endpackage

interface lwwreg_out_stream_if import lwwreg_pkg::*;;
    logic [3: 0] payload[2];
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface lwwreg_in_stream_if import lwwreg_pkg::*;;
    logic [3: 0] payload[2];
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module lwwreg import lwwreg_pkg::*;
 (
    input wire clk,
    input wire rst,
    lwwreg_out_stream_if.master out,
    lwwreg_in_stream_if.slave in
);
    // connect_rpc -exec amaranth-rpc yosys arq.LWWReg
    \arq.LWWReg  lwwreg_internal (
        .clk,
        .rst,
        .output__payload({<<4{out.p}}),
        .output__valid(out.valid),
        .output__ready(out.ready),
        .input__payload({<<4{in.p}}),
        .input__valid(in.valid)
    );

    assign in.ready = 1'd1;
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:250" *)
(* generator = "Amaranth" *)
module \arq.LWWReg (input__payload, input__valid, clk, rst, output__payload, output__valid, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$2 ;
  wire \$3 ;
  reg \$4 ;
  reg [7:0] \$5 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:252" *)
  reg [7:0] buffer = 8'h00;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:252" *)
  wire [3:0] \buffer[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:252" *)
  wire [3:0] \buffer[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:253" *)
  reg buffer_valid = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:244" *)
  input [7:0] input__payload;
  wire [7:0] input__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:244" *)
  wire [3:0] \input__payload[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:244" *)
  wire [3:0] \input__payload[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:244" *)
  output [7:0] output__payload;
  wire [7:0] output__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:244" *)
  wire [3:0] \output__payload[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:244" *)
  wire [3:0] \output__payload[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  assign \$3  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:261" *) \$2 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:253" *)
  always @(posedge clk)
    buffer_valid <= \$4 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:252" *)
  always @(posedge clk)
    buffer <= \$5 ;
  assign output__payload = input__valid ? (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:255" *) input__payload : buffer;
  assign output__valid = input__valid ? (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:256" *) input__valid : buffer_valid;
  assign \$1  = output__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:258" *) output__valid;
  assign \$2  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:261" *) output__ready;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$4  = buffer_valid;
    if (\$1 ) begin
      \$4  = 1'h0;
    end
    if (\$3 ) begin
      \$4  = 1'h1;
    end
    if (rst) begin
      \$4  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$5  = buffer;
    if (\$3 ) begin
      \$5  = input__payload;
    end
  end
  assign \output__payload[0]  = output__payload[3:0];
  assign \output__payload[1]  = output__payload[7:4];
  assign \input__payload[0]  = input__payload[3:0];
  assign \input__payload[1]  = input__payload[7:4];
  assign \buffer[0]  = buffer[3:0];
  assign \buffer[1]  = buffer[7:4];
endmodule


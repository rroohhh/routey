

package arq_receiver_pkg;
typedef struct packed {
    logic p;
    logic [1: 0] seq;
} arq_payload;

typedef struct packed {
    logic seq_is_valid;
    logic is_nack;
    logic [1: 0] seq;
} ack;
endpackage

interface arq_receiver_out_stream_if import arq_receiver_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_payload_stream_if import arq_receiver_pkg::*;;
    arq_payload payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_receiver_ack_if import arq_receiver_pkg::*;;
    ack p;
    logic trigger;
    logic did_trigger;

    modport master (
        output p,
        output trigger,
        input did_trigger
    );
    modport slave (
        input p,
        input trigger,
        output did_trigger
    );
    modport monitor (
        input p,
        input trigger,
        input did_trigger
    );
endinterface

module arq_receiver import arq_receiver_pkg::*;
 (
    input wire clk,
    input wire rst,
    input wire logic input_error,
    arq_receiver_out_stream_if.master out,
    arq_payload_stream_if.slave in,
    arq_receiver_ack_if.master ack
);
    // connect_rpc -exec amaranth-rpc yosys arq.ArqReceiver
    \arq.ArqReceiver  arq_receiver_internal (
        .clk,
        .rst,
        .input_error(input_error),
        .output__payload(out.p),
        .output__valid(out.valid),
        .output__ready(out.ready),
        .input__payload(in.p),
        .input__valid(in.valid),
        .input__ready(in.ready),
        .ack__p(ack.p),
        .ack__trigger(ack.trigger),
        .ack__did_trigger(ack.did_trigger)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post114, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:315" *)
(* generator = "Amaranth" *)
module \arq.ArqReceiver (output__ready, input__payload, input__valid, ack__did_trigger, clk, rst, output__payload, output__valid, input__ready, ack__p, ack__trigger, input_error);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire [2:0] \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire [2:0] \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  wire [1:0] \$22 ;
  wire [2:0] \$23 ;
  wire [3:0] \$24 ;
  wire \$25 ;
  wire \$26 ;
  wire \$27 ;
  wire \$28 ;
  wire \$29 ;
  wire \$3 ;
  wire \$30 ;
  reg \$31 ;
  reg [1:0] \$32 ;
  reg \$33 ;
  reg \$34 ;
  reg [1:0] \$35 ;
  reg \$36 ;
  wire \$4 ;
  wire \$5 ;
  wire \$6 ;
  wire [3:0] \$63 ;
  wire \$65 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:46" *)
  input ack__did_trigger;
  wire ack__did_trigger;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *)
  output [3:0] ack__p;
  wire [3:0] ack__p;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *)
  wire \ack__p.is_nack ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *)
  wire [1:0] \ack__p.seq ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *)
  wire \ack__p.seq_is_valid ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:45" *)
  output ack__trigger;
  reg ack__trigger = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:319" *)
  wire [1:0] expected_seq;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *)
  input [2:0] input__payload;
  wire [2:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *)
  wire \input__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *)
  wire [1:0] \input__payload.seq ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* annotation_text = "input error" *)
  (* debug_item = 32'd1 *)
  (* span_annotation = 32'd1 *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:308" *)
  input input_error;
  wire input_error;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:317" *)
  reg [1:0] last_seq = 2'h3;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:318" *)
  reg last_seq_valid = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:340" *)
  reg nack_scheduled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__payload;
  wire output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:209" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:369" *)
  reg [1:0] timeout_counter = 2'h0;
  (* annotation_text = "ack send timeout" *)
  (* debug_item = 32'd1 *)
  (* event_annotation = 32'd1 *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:417" *)
  wire timeout_occured;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:361" *)
  reg word_counter = 1'h0;
  assign \$1  = last_seq + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:320" *) 1'h1;
  assign \$2  = input__payload[1:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$1 [1:0];
  assign \$3  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$2 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:329" *) \$3 ;
  assign \$5  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:329" *) \$4 ;
  assign input__ready = output__ready | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:329" *) \$5 ;
  assign \$6  = input__payload[1:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$1 [1:0];
  assign output__valid = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$6 ;
  assign timeout_occured = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:418" *) timeout_counter;
  assign \$7  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:321" *) input__ready;
  assign \$8  = input__payload[1:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$1 [1:0];
  assign \$9  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$8 ;
  assign \$10  = \$7  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:324" *) \$9 ;
  assign \$11  = input__payload[1:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$1 [1:0];
  assign \$12  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$11 ;
  assign \$13  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:341" *) \$12 ;
  assign \$14  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:371" *) word_counter;
  assign \$15  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:374" *) timeout_counter;
  assign \$16  = timeout_counter - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:375" *) 1'h1;
  assign \$17  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:321" *) input__ready;
  assign \$18  = input__payload[1:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$1 [1:0];
  assign \$19  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$18 ;
  assign \$20  = \$17  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:380" *) \$19 ;
  assign \$22  = word_counter + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:387" *) 1'h1;
  assign \$23  = \$1 [1:0] - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:392" *) input__payload[1:0];
  wire [2:0] _0_ = $signed(\$23 ) % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:392" *) $signed(4'h4);
  assign \$63  = (\$23 [2] == 1'h0) || _0_ == 0 ? $signed(_0_) : $signed(4'h4) + $signed(_0_);
  assign \$25  = \$24 [2:0] > (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:392" *) 2'h2;
  assign \$26  = input__payload[1:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$1 [1:0];
  assign \$27  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:323" *) \$26 ;
  assign \$28  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:395" *) \$27 ;
  assign \$29  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:354" *) nack_scheduled;
  assign \$30  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:354" *) nack_scheduled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:318" *)
  always @(posedge clk)
    last_seq_valid <= \$31 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:317" *)
  always @(posedge clk)
    last_seq <= \$32 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:340" *)
  always @(posedge clk)
    nack_scheduled <= \$33 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:45" *)
  always @(posedge clk)
    ack__trigger <= \$34 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:369" *)
  always @(posedge clk)
    timeout_counter <= \$35 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:361" *)
  always @(posedge clk)
    word_counter <= \$36 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$31  = last_seq_valid;
    if (\$10 ) begin
      \$31  = 1'h1;
    end
    if (rst) begin
      \$31  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$32  = last_seq;
    if (\$10 ) begin
      \$32  = input__payload[1:0];
    end
    if (rst) begin
      \$32  = 2'h3;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$33  = nack_scheduled;
    if (\$13 ) begin
      \$33  = 1'h0;
    end
    if (input__valid) begin
      if (\$25 ) begin
        \$33  = 1'h1;
      end
    end
    if (input_error) begin
      \$33  = 1'h1;
    end
    if (rst) begin
      \$33  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$34  = 1'h0;
    (* full_case = 32'd1 *)
    if (\$14 ) begin
    end else begin
      (* full_case = 32'd1 *)
      if (\$15 ) begin
      end else begin
        \$34  = 1'h1;
      end
    end
    if (\$20 ) begin
      if (\$21 ) begin
        \$34  = 1'h1;
      end
    end
    if (input__valid) begin
      if (\$25 ) begin
        \$34  = \$29 ;
      end else if (\$28 ) begin
        \$34  = 1'h1;
      end
    end
    if (input_error) begin
      \$34  = \$30 ;
    end
    if (rst) begin
      \$34  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (\$14 ) begin
      \$35  = 2'h2;
    end else begin
      (* full_case = 32'd1 *)
      if (\$15 ) begin
        \$35  = \$16 [1:0];
      end else begin
        \$35  = 2'h2;
      end
    end
    if (\$20 ) begin
      if (\$21 ) begin
        \$35  = 2'h2;
      end
    end
    if (input__valid) begin
      if (\$25 ) begin
        \$35  = 2'h2;
      end else if (\$28 ) begin
        \$35  = 2'h2;
      end
    end
    if (ack__did_trigger) begin
      \$35  = 2'h2;
    end
    if (input_error) begin
      \$35  = 2'h2;
    end
    if (rst) begin
      \$35  = 2'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$36  = word_counter;
    (* full_case = 32'd1 *)
    if (\$14 ) begin
    end else begin
      (* full_case = 32'd1 *)
      if (\$15 ) begin
      end else begin
        \$36  = 1'h0;
      end
    end
    if (\$20 ) begin
      (* full_case = 32'd1 *)
      if (\$21 ) begin
        \$36  = 1'h0;
      end else begin
        \$36  = \$22 [0];
      end
    end
    if (ack__did_trigger) begin
      \$36  = 1'h0;
    end
    if (rst) begin
      \$36  = 1'h0;
    end
  end
  assign expected_seq = \$1 [1:0];
  assign output__payload = input__payload[2];
  assign \input__payload.seq  = input__payload[1:0];
  assign \input__payload.p  = input__payload[2];
  assign \ack__p.seq  = ack__p[1:0];
  assign \ack__p.is_nack  = ack__p[2];
  assign \ack__p.seq_is_valid  = ack__p[3];
  assign ack__p[2] = nack_scheduled;
  assign ack__p[3] = last_seq_valid;
  assign ack__p[1:0] = last_seq;
  assign \$21  = word_counter;
  assign \$65  = 1'h1;
  assign \$24  = \$63 ;
endmodule




package arq_sender_pkg;
typedef struct packed {
    logic p;
    logic [2: 0] seq;
} arq_payload;

typedef struct packed {
    logic seq_is_valid;
    logic is_nack;
    logic [2: 0] seq;
} ack;
endpackage

interface arq_sender_in_stream_if import arq_sender_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_payload_stream_if import arq_sender_pkg::*;;
    arq_payload payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface ack_stream_if import arq_sender_pkg::*;;
    ack payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module arq_sender import arq_sender_pkg::*;
 (
    input wire clk,
    input wire rst,
    arq_sender_in_stream_if.slave in,
    arq_payload_stream_if.master out,
    ack_stream_if.slave ack
);
    // connect_rpc -exec amaranth-rpc yosys arq.ArqSender
    \arq.ArqSender  arq_sender_internal (
        .clk,
        .rst,
        .input__payload(in.p),
        .input__valid(in.valid),
        .input__ready(in.ready),
        .output__payload(out.p),
        .output__valid(out.valid),
        .output__ready(out.ready),
        .ack__payload(ack.p),
        .ack__valid(ack.valid)
    );

    assign ack.ready = 1'd1;
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:60" *)
(* generator = "Amaranth" *)
module \arq.ArqSender (input__valid, output__ready, ack__payload, ack__valid, clk, rst, input__ready, output__payload, output__valid, input__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire [4:0] \$10 ;
  wire [4:0] \$101 ;
  wire \$103 ;
  wire \$11 ;
  wire [3:0] \$12 ;
  wire [3:0] \$13 ;
  wire [4:0] \$14 ;
  wire [4:0] \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire [3:0] \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  wire \$22 ;
  wire \$23 ;
  wire [4:0] \$24 ;
  wire \$25 ;
  wire \$26 ;
  wire [3:0] \$27 ;
  wire [3:0] \$28 ;
  wire [4:0] \$29 ;
  wire \$3 ;
  wire \$30 ;
  wire \$31 ;
  wire \$32 ;
  wire \$33 ;
  wire \$34 ;
  wire [3:0] \$35 ;
  wire [4:0] \$36 ;
  wire [4:0] \$37 ;
  wire \$38 ;
  wire \$39 ;
  wire \$4 ;
  reg [3:0] \$40 ;
  reg \$41 ;
  reg \$42 ;
  reg [2:0] \$43 ;
  reg [2:0] \$44 ;
  reg \$45 ;
  reg [2:0] \$46 ;
  reg [2:0] \$47 ;
  wire [3:0] \$5 ;
  wire \$6 ;
  wire [4:0] \$62 ;
  wire \$64 ;
  wire \$7 ;
  wire [4:0] \$71 ;
  wire \$73 ;
  wire \$8 ;
  wire [4:0] \$89 ;
  wire [3:0] \$9 ;
  wire \$91 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:53" *)
  input [4:0] ack__payload;
  wire [4:0] ack__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:53" *)
  wire \ack__payload.is_nack ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:53" *)
  wire [2:0] \ack__payload.seq ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:53" *)
  wire \ack__payload.seq_is_valid ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input ack__valid;
  wire ack__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:240" *)
  wire [1:0] buffer_read__addr;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:241" *)
  wire buffer_read__data;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:239" *)
  wire buffer_read__en;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:401" *)
  wire [1:0] buffer_write__addr;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:402" *)
  wire buffer_write__data;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:400" *)
  wire buffer_write__en;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:103" *)
  wire have_outstanding_to_send;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:402" *)
  input input__payload;
  wire input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* debug_item = 32'd1 *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:67" *)
  reg is_resend = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:120" *)
  reg last_was_empty_push = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:156" *)
  reg [2:0] next_read_ptr;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:65" *)
  reg [2:0] next_send_ptr;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:53" *)
  output [3:0] output__payload;
  wire [3:0] output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:53" *)
  wire \output__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:53" *)
  wire [2:0] \output__payload.seq ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:126" *)
  output output__valid;
  reg output__valid = 1'h0;
  (* capacity = 32'd4 *)
  (* debug_item = 32'd1 *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:194" *)
  wire [2:0] outstanding;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:76" *)
  wire pop;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:123" *)
  wire prefetch;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:74" *)
  wire push;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:63" *)
  reg [2:0] read_ptr = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:68" *)
  reg [2:0] resend_start = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* init = 1'h0 *)
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:126" *)
  wire send_outstanding;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:64" *)
  reg [2:0] send_ptr = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:121" *)
  reg send_ptr_moved;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:87" *)
  reg [3:0] timeout_counter = 4'h8;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:62" *)
  reg [2:0] write_ptr = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:70" *)
  reg [0:0] buffer [3:0];
  initial begin
    buffer[0] = 1'h0;
    buffer[1] = 1'h0;
    buffer[2] = 1'h0;
    buffer[3] = 1'h0;
  end
  always @(posedge clk) begin
    if (push)
      buffer[write_ptr[1:0]] <= input__payload;
  end
  reg [0:0] _0_;
  always @(posedge clk) begin
    if (prefetch) begin
      _0_ <= buffer[next_send_ptr[1:0]];
    end
  end
  assign buffer_read__data = _0_;
  assign \$36  = $signed(\$35 ) - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:183" *) $signed({ 1'h0, pop });
  wire [4:0] _1_ = $signed(\$36 ) % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:183" *) $signed(5'h08);
  assign \$101  = (\$36 [4] == 1'h0) || _1_ == 0 ? $signed(_1_) : $signed(5'h08) + $signed(_1_);
  assign \$38  = \$37 [3:0] <= (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:184" *) 3'h4;
  assign \$39  = next_read_ptr != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:164" *) write_ptr;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:87" *)
  always @(posedge clk)
    timeout_counter <= \$40 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:120" *)
  always @(posedge clk)
    last_was_empty_push <= \$41 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:126" *)
  always @(posedge clk)
    output__valid <= \$42 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:62" *)
  always @(posedge clk)
    write_ptr <= \$43 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:63" *)
  always @(posedge clk)
    read_ptr <= \$44 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:67" *)
  always @(posedge clk)
    is_resend <= \$45 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:68" *)
  always @(posedge clk)
    resend_start <= \$46 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:64" *)
  always @(posedge clk)
    send_ptr <= \$47 ;
  assign push = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:75" *) input__ready;
  assign pop = output__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:77" *) output__ready;
  assign have_outstanding_to_send = write_ptr != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:104" *) next_send_ptr;
  assign \$1  = write_ptr[2] != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:81" *) read_ptr[2];
  assign \$2  = write_ptr[1:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:81" *) read_ptr[1:0];
  assign \$3  = \$1  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:81" *) \$2 ;
  assign input__ready = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:113" *) \$3 ;
  assign \$4  = send_ptr_moved | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:124" *) last_was_empty_push;
  assign prefetch = \$4  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:124" *) have_outstanding_to_send;
  assign \$5  = send_ptr + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:154" *) 1'h1;
  assign \$6  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:88" *) timeout_counter;
  assign \$7  = next_read_ptr != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:164" *) write_ptr;
  assign \$9  = write_ptr - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:179" *) ack__payload[2:0];
  wire [3:0] _2_ = $signed(\$9 ) % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:179" *) $signed(5'h08);
  assign \$62  = (\$9 [3] == 1'h0) || _2_ == 0 ? $signed(_2_) : $signed(5'h08) + $signed(_2_);
  assign \$11  = \$10 [3:0] >= (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:179" *) 1'h1;
  assign \$12  = ack__payload[2:0] + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:180" *) \$11 ;
  assign \$13  = next_read_ptr - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:183" *) send_ptr;
  assign \$14  = $signed(\$13 ) - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:183" *) $signed({ 1'h0, pop });
  wire [4:0] _3_ = $signed(\$14 ) % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:183" *) $signed(5'h08);
  assign \$71  = (\$14 [4] == 1'h0) || _3_ == 0 ? $signed(_3_) : $signed(5'h08) + $signed(_3_);
  assign \$16  = \$15 [3:0] <= (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:184" *) 3'h4;
  assign \$17  = next_read_ptr != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:164" *) write_ptr;
  assign \$18  = write_ptr - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:197" *) read_ptr;
  assign \$19  = write_ptr == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:83" *) read_ptr;
  assign \$20  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:89" *) \$19 ;
  assign \$22  = \$21  | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:91" *) is_resend;
  assign \$23  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:94" *) timeout_counter;
  assign \$24  = timeout_counter - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:97" *) 1'h1;
  assign \$25  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:122" *) have_outstanding_to_send;
  assign \$26  = \$25  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:122" *) push;
  assign \$27  = write_ptr + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:151" *) 1'h1;
  assign \$28  = send_ptr - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:160" *) resend_start;
  wire [3:0] _4_ = $signed(\$28 ) % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:160" *) $signed(5'h08);
  assign \$89  = (\$28 [3] == 1'h0) || _4_ == 0 ? $signed(_4_) : $signed(5'h08) + $signed(_4_);
  assign \$30  = \$29 [3:0] < (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:160" *) 3'h4;
  assign \$31  = is_resend & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:160" *) \$30 ;
  assign \$32  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:88" *) timeout_counter;
  assign \$33  = next_read_ptr != (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:164" *) write_ptr;
  assign \$35  = next_read_ptr - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:183" *) send_ptr;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    next_send_ptr = send_ptr;
    if (pop) begin
      next_send_ptr = \$5 [2:0];
    end
    if (\$6 ) begin
      if (\$7 ) begin
        next_send_ptr = next_read_ptr;
      end
    end
    if (\$8 ) begin
      if (ack__payload[4]) begin
        if (\$16 ) begin
          next_send_ptr = next_read_ptr;
        end
      end
      if (ack__payload[3]) begin
        if (\$17 ) begin
          next_send_ptr = next_read_ptr;
        end
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    send_ptr_moved = 1'h0;
    if (pop) begin
      send_ptr_moved = 1'h1;
    end
    if (\$6 ) begin
      if (\$7 ) begin
        send_ptr_moved = 1'h1;
      end
    end
    if (\$8 ) begin
      if (ack__payload[4]) begin
        if (\$16 ) begin
          send_ptr_moved = 1'h1;
        end
      end
      if (ack__payload[3]) begin
        if (\$17 ) begin
          send_ptr_moved = 1'h1;
        end
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    next_read_ptr = read_ptr;
    if (\$8 ) begin
      if (ack__payload[4]) begin
        next_read_ptr = \$12 [2:0];
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (\$20 ) begin
      (* full_case = 32'd1 *)
      if (\$22 ) begin
        \$40  = 4'h8;
      end else begin
        (* full_case = 32'd1 *)
        if (\$23 ) begin
          \$40  = 4'h8;
        end else begin
          \$40  = \$24 [3:0];
        end
      end
    end else begin
      \$40  = 4'h8;
    end
    if (rst) begin
      \$40  = 4'h8;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$41  = \$26 ;
    if (rst) begin
      \$41  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$42  = output__valid;
    if (prefetch) begin
      \$42  = 1'h1;
    end
    if (pop) begin
      \$42  = prefetch;
    end
    if (\$32 ) begin
      if (\$33 ) begin
        \$42  = prefetch;
      end
    end
    if (\$34 ) begin
      if (ack__payload[4]) begin
        if (\$38 ) begin
          \$42  = prefetch;
        end
      end
      if (ack__payload[3]) begin
        if (\$39 ) begin
          \$42  = prefetch;
        end
      end
    end
    if (rst) begin
      \$42  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$43  = write_ptr;
    if (push) begin
      \$43  = \$27 [2:0];
    end
    if (rst) begin
      \$43  = 3'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$44  = next_read_ptr;
    if (rst) begin
      \$44  = 3'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$45  = is_resend;
    if (\$31 ) begin
      \$45  = 1'h0;
    end
    if (\$32 ) begin
      if (\$33 ) begin
        \$45  = 1'h1;
      end
    end
    if (\$34 ) begin
      if (ack__payload[3]) begin
        if (\$39 ) begin
          \$45  = 1'h1;
        end
      end
    end
    if (rst) begin
      \$45  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$46  = resend_start;
    if (\$32 ) begin
      if (\$33 ) begin
        \$46  = write_ptr;
      end
    end
    if (\$34 ) begin
      if (ack__payload[3]) begin
        if (\$39 ) begin
          \$46  = write_ptr;
        end
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$47  = next_send_ptr;
    if (rst) begin
      \$47  = 3'h0;
    end
  end
  assign buffer_write__en = push;
  assign buffer_write__addr = write_ptr[1:0];
  assign buffer_write__data = input__payload;
  assign buffer_read__en = prefetch;
  assign buffer_read__addr = next_send_ptr[1:0];
  assign send_outstanding = output__valid;
  assign outstanding = \$18 [2:0];
  assign \output__payload.seq  = output__payload[2:0];
  assign \output__payload.p  = output__payload[3];
  assign \ack__payload.seq  = ack__payload[2:0];
  assign \ack__payload.is_nack  = ack__payload[3];
  assign \ack__payload.seq_is_valid  = ack__payload[4];
  assign output__payload[2:0] = send_ptr;
  assign output__payload[3] = buffer_read__data;
  assign \$8  = ack__valid;
  assign \$64  = 1'h1;
  assign \$10  = \$62 ;
  assign \$73  = 1'h1;
  assign \$15  = \$71 ;
  assign \$21  = ack__valid;
  assign \$91  = 1'h1;
  assign \$29  = \$89 ;
  assign \$34  = ack__valid;
  assign \$103  = 1'h1;
  assign \$37  = \$101 ;
endmodule


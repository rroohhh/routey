

package arq_sender_pkg;
typedef struct packed {
    logic p;
    logic [3: 0] seq;
} arq_payload;

typedef struct packed {
    logic seq_is_valid;
    logic is_nack;
    logic [3: 0] seq;
} ack;
endpackage

interface arq_sender_in_stream_if import arq_sender_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_payload_stream_if import arq_sender_pkg::*;;
    arq_payload payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface ack_stream_if import arq_sender_pkg::*;;
    ack payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module arq_sender import arq_sender_pkg::*;
 (
    input wire clk,
    input wire rst,
    arq_sender_in_stream_if.slave in,
    arq_payload_stream_if.master out,
    ack_stream_if.slave ack
);
    // connect_rpc -exec amaranth-rpc yosys arq.ArqSender
    \arq.ArqSender  arq_sender_internal (
        .clk,
        .rst,
        .input__payload(in.p),
        .input__valid(in.valid),
        .input__ready(in.ready),
        .output__payload(out.p),
        .output__valid(out.valid),
        .output__ready(out.ready),
        .ack__payload(ack.p),
        .ack__valid(ack.valid)
    );

    assign ack.ready = 1'd1;
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:60" *)
(* generator = "Amaranth" *)
module \arq.ArqSender (input__valid, output__ready, ack__payload, ack__valid, clk, rst, input__ready, output__payload, output__valid, input__payload);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire \$17 ;
  wire \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire [4:0] \$20 ;
  wire \$21 ;
  wire \$22 ;
  wire \$23 ;
  wire \$24 ;
  wire \$25 ;
  wire \$26 ;
  wire \$27 ;
  wire \$28 ;
  wire \$29 ;
  wire \$3 ;
  wire \$30 ;
  wire \$31 ;
  wire \$32 ;
  wire \$33 ;
  wire \$34 ;
  wire [4:0] \$35 ;
  wire \$36 ;
  wire \$37 ;
  wire [4:0] \$38 ;
  wire [5:0] \$39 ;
  wire \$4 ;
  wire \$40 ;
  wire [4:0] \$41 ;
  wire [4:0] \$42 ;
  reg [4:0] \$43 ;
  reg \$44 ;
  reg \$45 ;
  reg [3:0] \$46 ;
  reg [3:0] \$47 ;
  reg \$48 ;
  reg [3:0] \$49 ;
  wire \$5 ;
  reg [3:0] \$50 ;
  wire [5:0] \$6 ;
  wire \$7 ;
  wire \$8 ;
  wire \$9 ;
  wire [5:0] \$92 ;
  wire \$94 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:53" *)
  input [5:0] ack__payload;
  wire [5:0] ack__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:53" *)
  wire \ack__payload.is_nack ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:53" *)
  wire [3:0] \ack__payload.seq ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:53" *)
  wire \ack__payload.seq_is_valid ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input ack__valid;
  wire ack__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:240" *)
  wire [2:0] buffer_read__addr;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:241" *)
  wire buffer_read__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:239" *)
  wire buffer_read__en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:401" *)
  wire [2:0] buffer_write__addr;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:402" *)
  wire buffer_write__data;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:400" *)
  wire buffer_write__en;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/memory.py:402" *)
  input input__payload;
  wire input__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* debug_item = 32'd1 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:67" *)
  reg is_resend = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:122" *)
  reg last_was_empty_push = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:121" *)
  reg nack;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:155" *)
  reg [3:0] next_read_ptr;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:65" *)
  reg [3:0] next_send_ptr;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:53" *)
  output [4:0] output__payload;
  wire [4:0] output__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:53" *)
  wire \output__payload.p ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:53" *)
  wire [3:0] \output__payload.seq ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:131" *)
  output output__valid;
  reg output__valid = 1'h0;
  (* capacity = 32'd8 *)
  (* debug_item = 32'd1 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:191" *)
  wire [3:0] outstanding;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:63" *)
  reg [3:0] read_ptr = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:68" *)
  reg [3:0] resend_start = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* init = 1'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:131" *)
  wire send_outstanding;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:64" *)
  reg [3:0] send_ptr = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:85" *)
  reg [4:0] timeout_counter = 5'h10;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:62" *)
  reg [3:0] write_ptr = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:70" *)
  reg [0:0] buffer [7:0];
  initial begin
    buffer[0] = 1'h0;
    buffer[1] = 1'h0;
    buffer[2] = 1'h0;
    buffer[3] = 1'h0;
    buffer[4] = 1'h0;
    buffer[5] = 1'h0;
    buffer[6] = 1'h0;
    buffer[7] = 1'h0;
  end
  always @(posedge clk) begin
    if (buffer_write__en)
      buffer[write_ptr[2:0]] <= input__payload;
  end
  reg [0:0] _0_;
  always @(posedge clk) begin
    if (buffer_read__en) begin
      _0_ <= buffer[next_send_ptr[2:0]];
    end
  end
  assign buffer_read__data = _0_;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:85" *)
  always @(posedge clk)
    timeout_counter <= \$43 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:122" *)
  always @(posedge clk)
    last_was_empty_push <= \$44 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:131" *)
  always @(posedge clk)
    output__valid <= \$45 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:62" *)
  always @(posedge clk)
    write_ptr <= \$46 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:63" *)
  always @(posedge clk)
    read_ptr <= \$47 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:67" *)
  always @(posedge clk)
    is_resend <= \$48 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:68" *)
  always @(posedge clk)
    resend_start <= \$49 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:64" *)
  always @(posedge clk)
    send_ptr <= \$50 ;
  assign \$1  = write_ptr == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:81" *) read_ptr;
  assign \$2  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:87" *) \$1 ;
  assign \$4  = \$3  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:89" *) is_resend;
  assign \$5  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:92" *) timeout_counter;
  assign \$6  = timeout_counter - (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:95" *) 1'h1;
  assign \$7  = write_ptr != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:101" *) next_send_ptr;
  assign \$8  = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:123" *) \$7 ;
  assign \$9  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:74" *) input__ready;
  assign \$10  = \$8  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:123" *) \$9 ;
  assign \$11  = output__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:75" *) output__ready;
  assign \$12  = \$11  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) nack;
  assign \$13  = \$12  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) last_was_empty_push;
  assign \$14  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:86" *) timeout_counter;
  assign \$15  = \$13  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) \$14 ;
  assign \$16  = write_ptr != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:101" *) next_send_ptr;
  assign \$17  = \$15  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) \$16 ;
  assign \$18  = output__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:75" *) output__ready;
  assign \$19  = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:74" *) input__ready;
  assign \$20  = write_ptr + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:150" *) 1'h1;
  assign \$21  = send_ptr == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:160" *) resend_start;
  assign \$22  = is_resend & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:160" *) \$21 ;
  assign \$23  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:86" *) timeout_counter;
  assign buffer_write__en = input__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:74" *) input__ready;
  assign \$25  = write_ptr[3] != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:79" *) read_ptr[3];
  assign \$26  = write_ptr[2:0] == (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:79" *) read_ptr[2:0];
  assign \$27  = \$25  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:79" *) \$26 ;
  assign input__ready = ~ (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:110" *) \$27 ;
  assign \$28  = output__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:75" *) output__ready;
  assign \$29  = \$28  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) nack;
  assign \$30  = \$29  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) last_was_empty_push;
  assign \$31  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:86" *) timeout_counter;
  assign \$32  = \$30  | (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) \$31 ;
  assign \$33  = write_ptr != (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:101" *) next_send_ptr;
  assign buffer_read__en = \$32  & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:124" *) \$33 ;
  assign \$34  = output__valid & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:75" *) output__ready;
  assign \$35  = send_ptr + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:153" *) 1'h1;
  assign \$36  = ! (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:86" *) timeout_counter;
  assign \$38  = write_ptr - (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:178" *) ack__payload[3:0];
  wire [4:0] _1_ = $signed(\$38 ) % (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:178" *) $signed(6'h10);
  assign \$92  = (\$38 [4] == 1'h0) || _1_ == 0 ? $signed(_1_) : $signed(6'h10) + $signed(_1_);
  assign \$40  = \$39 [4:0] > (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:178" *) 1'h1;
  assign \$41  = ack__payload[3:0] + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:179" *) \$40 ;
  assign \$42  = write_ptr - (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:194" *) read_ptr;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (\$2 ) begin
      (* full_case = 32'd1 *)
      if (\$4 ) begin
        \$43  = 5'h10;
      end else begin
        (* full_case = 32'd1 *)
        if (\$5 ) begin
          \$43  = 5'h10;
        end else begin
          \$43  = \$6 [4:0];
        end
      end
    end else begin
      \$43  = 5'h10;
    end
    if (rst) begin
      \$43  = 5'h10;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$44  = \$10 ;
    if (rst) begin
      \$44  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$45  = output__valid;
    if (\$17 ) begin
      \$45  = 1'h1;
    end else if (\$18 ) begin
      \$45  = 1'h0;
    end
    if (rst) begin
      \$45  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$46  = write_ptr;
    if (\$19 ) begin
      \$46  = \$20 [3:0];
    end
    if (rst) begin
      \$46  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$47  = next_read_ptr;
    if (rst) begin
      \$47  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$48  = is_resend;
    if (\$22 ) begin
      \$48  = 1'h0;
    end
    if (\$23 ) begin
      \$48  = 1'h1;
    end
    if (\$24 ) begin
      if (ack__payload[4]) begin
        \$48  = 1'h1;
      end
    end
    if (rst) begin
      \$48  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$49  = resend_start;
    if (\$23 ) begin
      \$49  = write_ptr;
    end
    if (\$24 ) begin
      if (ack__payload[4]) begin
        \$49  = write_ptr;
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$50  = next_send_ptr;
    if (rst) begin
      \$50  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    next_send_ptr = send_ptr;
    if (\$34 ) begin
      next_send_ptr = \$35 [3:0];
    end
    if (\$36 ) begin
      next_send_ptr = next_read_ptr;
    end
    if (\$37 ) begin
      if (ack__payload[4]) begin
        next_send_ptr = next_read_ptr;
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    next_read_ptr = read_ptr;
    if (\$37 ) begin
      if (ack__payload[5]) begin
        next_read_ptr = \$41 [3:0];
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    nack = 1'h0;
    if (\$37 ) begin
      if (ack__payload[4]) begin
        nack = 1'h1;
      end
    end
  end
  assign send_outstanding = output__valid;
  assign buffer_write__addr = write_ptr[2:0];
  assign buffer_write__data = input__payload;
  assign buffer_read__addr = next_send_ptr[2:0];
  assign outstanding = \$42 [3:0];
  assign \output__payload.seq  = output__payload[3:0];
  assign \output__payload.p  = output__payload[4];
  assign \ack__payload.seq  = ack__payload[3:0];
  assign \ack__payload.is_nack  = ack__payload[4];
  assign \ack__payload.seq_is_valid  = ack__payload[5];
  assign output__payload[3:0] = send_ptr;
  assign output__payload[4] = buffer_read__data;
  assign \$3  = ack__valid;
  assign \$24  = ack__valid;
  assign \$37  = ack__valid;
  assign \$94  = 1'h1;
  assign \$39  = \$92 ;
endmodule




package arq_receiver_pkg;
typedef struct packed {
    logic p;
    logic [2: 0] seq;
} arq_payload;

typedef struct packed {
    logic seq_is_valid;
    logic is_nack;
    logic [2: 0] seq;
} ack;
endpackage

interface arq_receiver_out_stream_if import arq_receiver_pkg::*;;
    logic payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_payload_stream_if import arq_receiver_pkg::*;;
    arq_payload payload;
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface arq_receiver_ack_if import arq_receiver_pkg::*;;
    ack p;
    logic trigger;
    logic did_trigger;

    modport master (
        output p,
        output trigger,
        input did_trigger
    );
    modport slave (
        input p,
        input trigger,
        output did_trigger
    );
    modport monitor (
        input p,
        input trigger,
        input did_trigger
    );
endinterface

module arq_receiver import arq_receiver_pkg::*;
 (
    input wire clk,
    input wire rst,
    input wire logic input_error,
    arq_receiver_out_stream_if.master out,
    arq_payload_stream_if.slave in,
    arq_receiver_ack_if.master ack
);
    // connect_rpc -exec amaranth-rpc yosys arq.ArqReceiver
    \arq.ArqReceiver  arq_receiver_internal (
        .clk,
        .rst,
        .input_error(input_error),
        .output__payload(out.p),
        .output__valid(out.valid),
        .output__ready(out.ready),
        .input__payload(in.p),
        .input__valid(in.valid),
        .input__ready(in.ready),
        .ack__p(ack.p),
        .ack__trigger(ack.trigger),
        .ack__did_trigger(ack.did_trigger)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:301" *)
(* generator = "Amaranth" *)
module \arq.ArqReceiver (output__ready, input__payload, input__valid, ack__did_trigger, clk, rst, output__payload, output__valid, input__ready, ack__p, ack__trigger, input_error);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire [3:0] \$1 ;
  wire \$10 ;
  wire \$11 ;
  wire \$12 ;
  wire \$13 ;
  wire \$14 ;
  wire \$15 ;
  wire \$16 ;
  wire [3:0] \$17 ;
  wire [4:0] \$18 ;
  wire \$19 ;
  wire \$2 ;
  wire \$20 ;
  wire \$21 ;
  wire \$22 ;
  wire \$23 ;
  wire \$24 ;
  wire \$25 ;
  wire \$26 ;
  wire \$27 ;
  wire \$28 ;
  wire \$29 ;
  wire \$3 ;
  wire \$30 ;
  wire [3:0] \$31 ;
  wire \$32 ;
  wire \$33 ;
  wire \$34 ;
  wire \$35 ;
  wire \$36 ;
  wire [1:0] \$37 ;
  wire [3:0] \$38 ;
  wire [4:0] \$39 ;
  wire \$4 ;
  wire \$40 ;
  wire \$41 ;
  wire \$42 ;
  wire \$43 ;
  reg \$44 ;
  reg [2:0] \$45 ;
  reg \$46 ;
  reg [2:0] \$47 ;
  reg \$48 ;
  wire \$5 ;
  wire \$6 ;
  wire [4:0] \$68 ;
  wire \$7 ;
  wire \$70 ;
  wire \$8 ;
  wire \$9 ;
  wire [4:0] \$93 ;
  wire \$95 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:46" *)
  input ack__did_trigger;
  wire ack__did_trigger;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:293" *)
  output [4:0] ack__p;
  reg [4:0] ack__p;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:293" *)
  wire \ack__p.is_nack ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:293" *)
  wire [2:0] \ack__p.seq ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:293" *)
  wire \ack__p.seq_is_valid ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:45" *)
  output ack__trigger;
  reg ack__trigger;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:305" *)
  wire [2:0] expected_seq;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:293" *)
  input [3:0] input__payload;
  wire [3:0] input__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:293" *)
  wire \input__payload.p ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:293" *)
  wire [2:0] \input__payload.seq ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  output input__ready;
  wire input__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:294" *)
  input input_error;
  wire input_error;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:303" *)
  reg [2:0] last_seq = 3'h7;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:304" *)
  reg last_seq_valid = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:326" *)
  reg nack_scheduled = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:327" *)
  reg next_nack_scheduled;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:48" *)
  output output__payload;
  wire output__payload;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  output output__valid;
  wire output__valid;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:357" *)
  reg [2:0] timeout_counter = 3'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:349" *)
  reg word_counter = 1'h0;
  assign \$42  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$41 ;
  assign \$43  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:383" *) \$42 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:304" *)
  always @(posedge clk)
    last_seq_valid <= \$44 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:303" *)
  always @(posedge clk)
    last_seq <= \$45 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:326" *)
  always @(posedge clk)
    nack_scheduled <= \$46 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:357" *)
  always @(posedge clk)
    timeout_counter <= \$47 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:349" *)
  always @(posedge clk)
    word_counter <= \$48 ;
  assign \$1  = last_seq + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:306" *) 1'h1;
  assign \$2  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  assign \$3  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$2 ;
  assign \$4  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:315" *) \$3 ;
  assign \$5  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:315" *) \$4 ;
  assign input__ready = output__ready | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:315" *) \$5 ;
  assign \$6  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  assign output__valid = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$6 ;
  assign \$7  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  assign \$8  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$7 ;
  assign \$9  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:330" *) \$8 ;
  assign \$10  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:359" *) word_counter;
  assign \$11  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:362" *) timeout_counter;
  assign \$12  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *) input__ready;
  assign \$13  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  assign \$14  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$13 ;
  assign \$15  = \$12  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:368" *) \$14 ;
  assign \$17  = \$1 [2:0] - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:380" *) input__payload[2:0];
  wire [3:0] _0_ = $signed(\$17 ) % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:380" *) $signed(5'h08);
  assign \$68  = (\$17 [3] == 1'h0) || _0_ == 0 ? $signed(_0_) : $signed(5'h08) + $signed(_0_);
  assign \$19  = \$18 [3:0] > (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:380" *) 3'h4;
  assign \$20  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  assign \$21  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$20 ;
  assign \$22  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:383" *) \$21 ;
  assign \$23  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:342" *) nack_scheduled;
  assign \$24  = ~ (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:342" *) nack_scheduled;
  assign \$25  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *) input__ready;
  assign \$26  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  assign \$27  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$26 ;
  assign \$28  = \$25  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:310" *) \$27 ;
  assign \$29  = ! (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:359" *) word_counter;
  assign \$30  = | (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:362" *) timeout_counter;
  assign \$31  = timeout_counter - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:363" *) 1'h1;
  assign \$32  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:307" *) input__ready;
  assign \$33  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  assign \$34  = input__valid & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$33 ;
  assign \$35  = \$32  & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:368" *) \$34 ;
  assign \$37  = word_counter + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:375" *) 1'h1;
  assign \$38  = \$1 [2:0] - (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:380" *) input__payload[2:0];
  wire [3:0] _1_ = $signed(\$38 ) % (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:380" *) $signed(5'h08);
  assign \$93  = (\$38 [3] == 1'h0) || _1_ == 0 ? $signed(_1_) : $signed(5'h08) + $signed(_1_);
  assign \$40  = \$39 [3:0] > (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:380" *) 3'h4;
  assign \$41  = input__payload[2:0] == (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:309" *) \$1 [2:0];
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    ack__p[2:0] = last_seq;
    if (\$15 ) begin
      if (\$16 ) begin
        ack__p[2:0] = \$1 [2:0];
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    next_nack_scheduled = nack_scheduled;
    if (\$9 ) begin
      next_nack_scheduled = 1'h0;
    end
    if (input__valid) begin
      if (\$19 ) begin
        next_nack_scheduled = 1'h1;
      end
    end
    if (input_error) begin
      next_nack_scheduled = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    ack__trigger = 1'h0;
    (* full_case = 32'd1 *)
    if (\$10 ) begin
    end else begin
      (* full_case = 32'd1 *)
      if (\$11 ) begin
      end else begin
        ack__trigger = 1'h1;
      end
    end
    if (\$15 ) begin
      if (\$16 ) begin
        ack__trigger = 1'h1;
      end
    end
    if (input__valid) begin
      if (\$19 ) begin
        ack__trigger = \$23 ;
      end else if (\$22 ) begin
        ack__trigger = 1'h1;
      end
    end
    if (input_error) begin
      ack__trigger = \$24 ;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$44  = last_seq_valid;
    if (\$28 ) begin
      \$44  = 1'h1;
    end
    if (rst) begin
      \$44  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$45  = last_seq;
    if (\$28 ) begin
      \$45  = input__payload[2:0];
    end
    if (rst) begin
      \$45  = 3'h7;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$46  = next_nack_scheduled;
    if (rst) begin
      \$46  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (\$29 ) begin
      \$47  = 3'h4;
    end else begin
      (* full_case = 32'd1 *)
      if (\$30 ) begin
        \$47  = \$31 [2:0];
      end else begin
        \$47  = 3'h4;
      end
    end
    if (\$35 ) begin
      if (\$36 ) begin
        \$47  = 3'h4;
      end
    end
    if (input__valid) begin
      if (\$40 ) begin
        \$47  = 3'h4;
      end else if (\$43 ) begin
        \$47  = 3'h4;
      end
    end
    if (ack__did_trigger) begin
      \$47  = 3'h4;
    end
    if (input_error) begin
      \$47  = 3'h4;
    end
    if (rst) begin
      \$47  = 3'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$48  = word_counter;
    (* full_case = 32'd1 *)
    if (\$29 ) begin
    end else begin
      (* full_case = 32'd1 *)
      if (\$30 ) begin
      end else begin
        \$48  = 1'h0;
      end
    end
    if (\$35 ) begin
      (* full_case = 32'd1 *)
      if (\$36 ) begin
        \$48  = 1'h0;
      end else begin
        \$48  = \$37 [0];
      end
    end
    if (ack__did_trigger) begin
      \$48  = 1'h0;
    end
    if (rst) begin
      \$48  = 1'h0;
    end
  end
  assign expected_seq = \$1 [2:0];
  assign output__payload = input__payload[3];
  assign \input__payload.seq  = input__payload[2:0];
  assign \input__payload.p  = input__payload[3];
  assign \ack__p.seq  = ack__p[2:0];
  assign \ack__p.is_nack  = ack__p[3];
  assign \ack__p.seq_is_valid  = ack__p[4];
  always @*
    ack__p[3] = next_nack_scheduled;
  always @*
    ack__p[4] = last_seq_valid;
  assign \$16  = word_counter;
  assign \$70  = 1'h1;
  assign \$18  = \$68 ;
  assign \$36  = word_counter;
  assign \$95  = 1'h1;
  assign \$39  = \$93 ;
endmodule


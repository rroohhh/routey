

package multi_queue_credit_counter_rx_pkg;
typedef struct packed {
    logic ready;
    logic valid;
} stream_monitor;
endpackage

interface multi_queue_credit_counter_rx_credit_out_if import multi_queue_credit_counter_rx_pkg::*;;
    logic [3: 0] credit[2];
    logic did_trigger;
    logic trigger;

    modport master (
        output credit,
        input did_trigger,
        output trigger
    );
    modport slave (
        input credit,
        output did_trigger,
        input trigger
    );
    modport monitor (
        input credit,
        input did_trigger,
        input trigger
    );
endinterface

module multi_queue_credit_counter_rx import multi_queue_credit_counter_rx_pkg::*;
 (
    input wire clk,
    input wire rst,
    input wire stream_monitor fifo_output_monitor[2],
    multi_queue_credit_counter_rx_credit_out_if.master credit_out
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueCreditCounterRX
    \arq.MultiQueueCreditCounterRX  multi_queue_credit_counter_rx_internal (
        .clk,
        .rst,
        .fifo_output_monitor__0(fifo_output_monitor[0]),
        .fifo_output_monitor__1(fifo_output_monitor[1]),
        .credit_out__credit({<<4{credit_out.credit}}),
        .credit_out__did_trigger(credit_out.did_trigger),
        .credit_out__trigger(credit_out.trigger)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:865" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueCreditCounterRX (fifo_output_monitor__1, credit_out__did_trigger, clk, rst, credit_out__credit, credit_out__trigger, fifo_output_monitor__0);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  reg [3:0] \$10 ;
  reg [3:0] \$11 ;
  reg \$12 ;
  wire \$2 ;
  wire \$3 ;
  wire \$4 ;
  wire [4:0] \$5 ;
  wire \$6 ;
  wire [4:0] \$7 ;
  wire \$8 ;
  wire [1:0] \$9 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *)
  output [7:0] credit_out__credit;
  wire [7:0] credit_out__credit;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *)
  wire [3:0] \credit_out__credit[0] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:856" *)
  wire [3:0] \credit_out__credit[1] ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:849" *)
  input credit_out__did_trigger;
  wire credit_out__did_trigger;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:850" *)
  output credit_out__trigger;
  reg credit_out__trigger;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:877" *)
  reg credit_trigger_timer = 1'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:868" *)
  reg did_read;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  input [1:0] fifo_output_monitor__0;
  wire [1:0] fifo_output_monitor__0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__0.ready ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__0.valid ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  input [1:0] fifo_output_monitor__1;
  wire [1:0] fifo_output_monitor__1;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__1.ready ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__1.valid ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:867" *)
  reg [3:0] read_ptr_0 = 4'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:867" *)
  reg [3:0] read_ptr_1 = 4'h0;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  assign \$1  = fifo_output_monitor__0[0] & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:872" *) fifo_output_monitor__0[1];
  assign \$2  = fifo_output_monitor__1[0] & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:872" *) fifo_output_monitor__1[1];
  assign \$4  = fifo_output_monitor__0[0] & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:872" *) fifo_output_monitor__0[1];
  assign \$5  = read_ptr_0 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:873" *) 1'h1;
  assign \$6  = fifo_output_monitor__1[0] & (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:872" *) fifo_output_monitor__1[1];
  assign \$7  = read_ptr_1 + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:873" *) 1'h1;
  assign \$9  = credit_trigger_timer + (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:886" *) did_read;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:867" *)
  always @(posedge clk)
    read_ptr_0 <= \$10 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:867" *)
  always @(posedge clk)
    read_ptr_1 <= \$11 ;
  (* src = "/data/study/master/thesis/work/toplevel_xcelium/fatmeshy/units/config_router/arq.py:877" *)
  always @(posedge clk)
    credit_trigger_timer <= \$12 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    did_read = 1'h0;
    if (\$1 ) begin
      did_read = 1'h1;
    end
    if (\$2 ) begin
      did_read = 1'h1;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    credit_out__trigger = 1'h0;
    (* full_case = 32'd1 *)
    if (credit_out__did_trigger) begin
    end else begin
      if (\$3 ) begin
        credit_out__trigger = 1'h1;
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$10  = read_ptr_0;
    if (\$4 ) begin
      \$10  = \$5 [3:0];
    end
    if (rst) begin
      \$10  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$11  = read_ptr_1;
    if (\$6 ) begin
      \$11  = \$7 [3:0];
    end
    if (rst) begin
      \$11  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (credit_out__did_trigger) begin
      \$12  = 1'h0;
    end else begin
      (* full_case = 32'd1 *)
      if (\$8 ) begin
        \$12  = 1'h0;
      end else begin
        \$12  = \$9 [0];
      end
    end
    if (rst) begin
      \$12  = 1'h0;
    end
  end
  assign \fifo_output_monitor__0.valid  = fifo_output_monitor__0[0];
  assign \fifo_output_monitor__0.ready  = fifo_output_monitor__0[1];
  assign \fifo_output_monitor__1.valid  = fifo_output_monitor__1[0];
  assign \fifo_output_monitor__1.ready  = fifo_output_monitor__1[1];
  assign \credit_out__credit[0]  = credit_out__credit[3:0];
  assign \credit_out__credit[1]  = credit_out__credit[7:4];
  assign credit_out__credit[7:4] = read_ptr_1;
  assign credit_out__credit[3:0] = read_ptr_0;
  assign \$3  = credit_trigger_timer;
  assign \$8  = credit_trigger_timer;
endmodule


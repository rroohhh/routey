

package lwwreg_pkg;

endpackage

interface lwwreg_out_stream_if import lwwreg_pkg::*;;
    logic [3: 0] payload[2];
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

interface lwwreg_in_stream_if import lwwreg_pkg::*;;
    logic [3: 0] payload[2];
    logic valid;
    logic ready;

    modport master (
        output .p(payload),
        output valid,
        input ready
    );
    modport slave (
        input .p(payload),
        input valid,
        output ready
    );
    modport monitor (
        input .p(payload),
        input valid,
        input ready
    );
endinterface

module lwwreg import lwwreg_pkg::*;
 (
    input wire clk,
    input wire rst,
    lwwreg_out_stream_if.master out,
    output wire logic buffer_valid,
    lwwreg_in_stream_if.slave in
);
    // connect_rpc -exec amaranth-rpc yosys arq.LWWReg
    \arq.LWWReg  lwwreg_internal (
        .clk,
        .rst,
        .output__payload({<<4{out.p}}),
        .output__valid(out.valid),
        .output__ready(out.ready),
        .buffer_valid(buffer_valid),
        .input__payload({<<4{in.p}}),
        .input__valid(in.valid)
    );

    assign in.ready = 1'd1;
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:267" *)
(* generator = "Amaranth" *)
module \arq.LWWReg (input__payload, input__valid, clk, rst, output__payload, output__valid, buffer_valid, output__ready);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  wire \$2 ;
  reg \$3 ;
  reg [7:0] \$4 ;
  (* init = 8'h00 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:269" *)
  wire [7:0] buffer;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:269" *)
  wire [3:0] \buffer[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:269" *)
  wire [3:0] \buffer[1] ;
  (* init = 1'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:262" *)
  output buffer_valid;
  wire buffer_valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:260" *)
  input [7:0] input__payload;
  wire [7:0] input__payload;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:260" *)
  wire [3:0] \input__payload[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:260" *)
  wire [3:0] \input__payload[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:49" *)
  input input__valid;
  wire input__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:269" *)
  output [7:0] output__payload;
  reg [7:0] output__payload = 8'h00;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:260" *)
  wire [3:0] \output__payload[0] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:260" *)
  wire [3:0] \output__payload[1] ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/stream.py:50" *)
  input output__ready;
  wire output__ready;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:262" *)
  output output__valid;
  reg output__valid = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:269" *)
  always @(posedge clk)
    output__payload <= \$4 ;
  assign \$1  = output__ready & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:275" *) output__valid;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:262" *)
  always @(posedge clk)
    output__valid <= \$3 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$3  = output__valid;
    if (\$1 ) begin
      \$3  = 1'h0;
    end
    if (\$2 ) begin
      \$3  = 1'h1;
    end
    if (rst) begin
      \$3  = 1'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$4  = output__payload;
    if (\$2 ) begin
      \$4  = input__payload;
    end
  end
  assign buffer = output__payload;
  assign buffer_valid = output__valid;
  assign \output__payload[0]  = output__payload[3:0];
  assign \output__payload[1]  = output__payload[7:4];
  assign \input__payload[0]  = input__payload[3:0];
  assign \input__payload[1]  = input__payload[7:4];
  assign \buffer[0]  = output__payload[3:0];
  assign \buffer[1]  = output__payload[7:4];
  assign \$2  = input__valid;
endmodule




package multi_queue_credit_counter_rx_pkg;
typedef struct packed {
    logic ready;
    logic valid;
    logic p;
} stream_monitor;
endpackage

module multi_queue_credit_counter_rx import multi_queue_credit_counter_rx_pkg::*;
 (
    input wire clk,
    input wire rst,
    input wire stream_monitor fifo_output_monitor[2],
    output wire logic [3: 0] credit_out[2],
    input wire logic credit_out_did_trigger,
    output wire logic credit_out_trigger
);
    // connect_rpc -exec amaranth-rpc yosys arq.MultiQueueCreditCounterRX
    \arq.MultiQueueCreditCounterRX  multi_queue_credit_counter_rx_internal (
        .clk,
        .rst,
        .fifo_output_monitor__0(fifo_output_monitor[0]),
        .fifo_output_monitor__1(fifo_output_monitor[1]),
        .credit_out__0(credit_out[0]),
        .credit_out__1(credit_out[1]),
        .credit_out_did_trigger(credit_out_did_trigger),
        .credit_out_trigger(credit_out_trigger)
    );
endmodule
/* Generated by Amaranth Yosys 0.50 (PyPI ver 0.50.0.0.post108, git sha1 b5170e139) */

(* top =  1  *)
(* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:795" *)
(* generator = "Amaranth" *)
module \arq.MultiQueueCreditCounterRX (fifo_output_monitor__1, credit_out_did_trigger, clk, rst, credit_out__0, credit_out__1, credit_out_trigger, fifo_output_monitor__0);
  reg \$auto$verilog_backend.cc:2355:dump_module$1  = 0;
  wire \$1 ;
  reg \$10 ;
  wire \$2 ;
  wire [4:0] \$3 ;
  wire \$4 ;
  wire [4:0] \$5 ;
  wire \$6 ;
  wire [1:0] \$7 ;
  reg [3:0] \$8 ;
  reg [3:0] \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input clk;
  wire clk;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:797" *)
  output [3:0] credit_out__0;
  reg [3:0] credit_out__0 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:797" *)
  output [3:0] credit_out__1;
  reg [3:0] credit_out__1 = 4'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:787" *)
  input credit_out_did_trigger;
  wire credit_out_did_trigger;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:788" *)
  output credit_out_trigger;
  reg credit_out_trigger;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:805" *)
  reg credit_trigger_timer = 1'h0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  input [2:0] fifo_output_monitor__0;
  wire [2:0] fifo_output_monitor__0;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__0.p ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__0.ready ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__0.valid ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  input [2:0] fifo_output_monitor__1;
  wire [2:0] fifo_output_monitor__1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__1.p ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__1.ready ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/lib/wiring.py:1695" *)
  wire \fifo_output_monitor__1.valid ;
  (* init = 4'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:797" *)
  wire [3:0] read_ptr_0;
  (* init = 4'h0 *)
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:797" *)
  wire [3:0] read_ptr_1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/.venv/lib64/python3.9/site-packages/amaranth/hdl/_ir.py:211" *)
  input rst;
  wire rst;
  assign \$2  = fifo_output_monitor__0[1] & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:801" *) fifo_output_monitor__0[2];
  assign \$3  = credit_out__0 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:802" *) 1'h1;
  assign \$4  = fifo_output_monitor__1[1] & (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:801" *) fifo_output_monitor__1[2];
  assign \$5  = credit_out__1 + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:802" *) 1'h1;
  assign \$7  = credit_trigger_timer + (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:814" *) 1'h1;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:797" *)
  always @(posedge clk)
    credit_out__0 <= \$8 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:797" *)
  always @(posedge clk)
    credit_out__1 <= \$9 ;
  (* src = "/hyperfast/home/rheinema/master/fatmeshy/units/config_router/arq.py:805" *)
  always @(posedge clk)
    credit_trigger_timer <= \$10 ;
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    credit_out_trigger = 1'h0;
    (* full_case = 32'd1 *)
    if (credit_out_did_trigger) begin
    end else begin
      if (\$1 ) begin
        credit_out_trigger = 1'h1;
      end
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$8  = credit_out__0;
    if (\$2 ) begin
      \$8  = \$3 [3:0];
    end
    if (rst) begin
      \$8  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    \$9  = credit_out__1;
    if (\$4 ) begin
      \$9  = \$5 [3:0];
    end
    if (rst) begin
      \$9  = 4'h0;
    end
  end
  always @* begin
    if (\$auto$verilog_backend.cc:2355:dump_module$1 ) begin end
    (* full_case = 32'd1 *)
    if (credit_out_did_trigger) begin
      \$10  = 1'h0;
    end else begin
      (* full_case = 32'd1 *)
      if (\$6 ) begin
        \$10  = 1'h0;
      end else begin
        \$10  = \$7 [0];
      end
    end
    if (rst) begin
      \$10  = 1'h0;
    end
  end
  assign read_ptr_0 = credit_out__0;
  assign read_ptr_1 = credit_out__1;
  assign \fifo_output_monitor__0.p  = fifo_output_monitor__0[0];
  assign \fifo_output_monitor__0.valid  = fifo_output_monitor__0[1];
  assign \fifo_output_monitor__0.ready  = fifo_output_monitor__0[2];
  assign \fifo_output_monitor__1.p  = fifo_output_monitor__1[0];
  assign \fifo_output_monitor__1.valid  = fifo_output_monitor__1[1];
  assign \fifo_output_monitor__1.ready  = fifo_output_monitor__1[2];
  assign \$1  = credit_trigger_timer;
  assign \$6  = credit_trigger_timer;
endmodule

